//Generate the verilog at 2025-07-28T18:07:49 by iSTA.
module ysyx_25040111 (
clock,
reset
);

input clock ;
input reset ;




endmodule
