//Generate the verilog at 2025-10-20T11:01:39 by iSTA.
module ysyx_25040111 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire de_ard_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire ea_err ;
wire ea_rsign ;
wire exe_valid ;
wire exu_valid ;
wire flush_$_OR__Y_B ;
wire icah_valid ;
wire idu_ready ;
wire ifu_ready ;
wire io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_B ;
wire io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_B ;
wire io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_B ;
wire io_master_araddr_$_NOT__Y_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_A_$_MUX__Y_B ;
wire io_master_bvalid_$_OR__B_Y ;
wire io_master_rready_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A ;
wire io_master_rready_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_MUX__Y_B ;
wire \u_arbiter.rsign ;
wire \u_arbiter.rvalid ;
wire \u_arbiter.rvalid_$_SDFFE_PP0P__Q_E ;
wire \u_arbiter.working ;
wire \u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ;
wire \u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_AND__A_Y ;
wire \u_arbiter.working_$_SDFFE_PP0P__Q_E ;
wire \u_arbiter.wvalid ;
wire \u_arbiter.wvalid_$_SDFFE_PP0P__Q_E ;
wire \u_csr.csr[0][0] ;
wire \u_csr.csr[0][10] ;
wire \u_csr.csr[0][11] ;
wire \u_csr.csr[0][12] ;
wire \u_csr.csr[0][13] ;
wire \u_csr.csr[0][14] ;
wire \u_csr.csr[0][15] ;
wire \u_csr.csr[0][16] ;
wire \u_csr.csr[0][17] ;
wire \u_csr.csr[0][18] ;
wire \u_csr.csr[0][19] ;
wire \u_csr.csr[0][1] ;
wire \u_csr.csr[0][20] ;
wire \u_csr.csr[0][21] ;
wire \u_csr.csr[0][22] ;
wire \u_csr.csr[0][23] ;
wire \u_csr.csr[0][24] ;
wire \u_csr.csr[0][25] ;
wire \u_csr.csr[0][26] ;
wire \u_csr.csr[0][27] ;
wire \u_csr.csr[0][28] ;
wire \u_csr.csr[0][29] ;
wire \u_csr.csr[0][2] ;
wire \u_csr.csr[0][30] ;
wire \u_csr.csr[0][31] ;
wire \u_csr.csr[0][3] ;
wire \u_csr.csr[0][4] ;
wire \u_csr.csr[0][5] ;
wire \u_csr.csr[0][6] ;
wire \u_csr.csr[0][7] ;
wire \u_csr.csr[0][8] ;
wire \u_csr.csr[0][9] ;
wire \u_csr.csr[1][0] ;
wire \u_csr.csr[1][10] ;
wire \u_csr.csr[1][11] ;
wire \u_csr.csr[1][12] ;
wire \u_csr.csr[1][13] ;
wire \u_csr.csr[1][14] ;
wire \u_csr.csr[1][15] ;
wire \u_csr.csr[1][16] ;
wire \u_csr.csr[1][17] ;
wire \u_csr.csr[1][18] ;
wire \u_csr.csr[1][19] ;
wire \u_csr.csr[1][1] ;
wire \u_csr.csr[1][20] ;
wire \u_csr.csr[1][21] ;
wire \u_csr.csr[1][22] ;
wire \u_csr.csr[1][23] ;
wire \u_csr.csr[1][24] ;
wire \u_csr.csr[1][25] ;
wire \u_csr.csr[1][26] ;
wire \u_csr.csr[1][27] ;
wire \u_csr.csr[1][28] ;
wire \u_csr.csr[1][29] ;
wire \u_csr.csr[1][2] ;
wire \u_csr.csr[1][30] ;
wire \u_csr.csr[1][31] ;
wire \u_csr.csr[1][3] ;
wire \u_csr.csr[1][4] ;
wire \u_csr.csr[1][5] ;
wire \u_csr.csr[1][6] ;
wire \u_csr.csr[1][7] ;
wire \u_csr.csr[1][8] ;
wire \u_csr.csr[1][9] ;
wire \u_csr.csr[2][0] ;
wire \u_csr.csr[2][10] ;
wire \u_csr.csr[2][11] ;
wire \u_csr.csr[2][12] ;
wire \u_csr.csr[2][13] ;
wire \u_csr.csr[2][14] ;
wire \u_csr.csr[2][15] ;
wire \u_csr.csr[2][16] ;
wire \u_csr.csr[2][17] ;
wire \u_csr.csr[2][18] ;
wire \u_csr.csr[2][19] ;
wire \u_csr.csr[2][1] ;
wire \u_csr.csr[2][20] ;
wire \u_csr.csr[2][21] ;
wire \u_csr.csr[2][22] ;
wire \u_csr.csr[2][23] ;
wire \u_csr.csr[2][24] ;
wire \u_csr.csr[2][25] ;
wire \u_csr.csr[2][26] ;
wire \u_csr.csr[2][27] ;
wire \u_csr.csr[2][28] ;
wire \u_csr.csr[2][29] ;
wire \u_csr.csr[2][2] ;
wire \u_csr.csr[2][30] ;
wire \u_csr.csr[2][31] ;
wire \u_csr.csr[2][3] ;
wire \u_csr.csr[2][4] ;
wire \u_csr.csr[2][5] ;
wire \u_csr.csr[2][6] ;
wire \u_csr.csr[2][7] ;
wire \u_csr.csr[2][8] ;
wire \u_csr.csr[2][9] ;
wire \u_csr.csr[3][0] ;
wire \u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y ;
wire \u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_exu.alu_p2_$_SDFFE_PP0P__Q_E ;
wire \u_exu.exe_end_$_ANDNOT__B_Y ;
wire \u_exu.exe_end_$_SDFFE_PP0P__Q_E ;
wire \u_exu.exe_start ;
wire \u_exu.exe_start_$_SDFFE_PP0P__Q_E ;
wire \u_exu.jmpc_ok ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_1_B ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_B ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ;
wire \u_exu.opt_$_NOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B ;
wire \u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ;
wire \u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ;
wire \u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B_$_MUX__B_A_$_NAND__Y_B ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_Y_$_MUX__B_A_$_NOR__Y_A_$_ANDNOT__Y_B ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_icache.cblocks[0][0] ;
wire \u_icache.cblocks[0][10] ;
wire \u_icache.cblocks[0][11] ;
wire \u_icache.cblocks[0][12] ;
wire \u_icache.cblocks[0][13] ;
wire \u_icache.cblocks[0][14] ;
wire \u_icache.cblocks[0][15] ;
wire \u_icache.cblocks[0][16] ;
wire \u_icache.cblocks[0][17] ;
wire \u_icache.cblocks[0][18] ;
wire \u_icache.cblocks[0][19] ;
wire \u_icache.cblocks[0][1] ;
wire \u_icache.cblocks[0][20] ;
wire \u_icache.cblocks[0][21] ;
wire \u_icache.cblocks[0][22] ;
wire \u_icache.cblocks[0][23] ;
wire \u_icache.cblocks[0][24] ;
wire \u_icache.cblocks[0][25] ;
wire \u_icache.cblocks[0][26] ;
wire \u_icache.cblocks[0][27] ;
wire \u_icache.cblocks[0][28] ;
wire \u_icache.cblocks[0][29] ;
wire \u_icache.cblocks[0][2] ;
wire \u_icache.cblocks[0][30] ;
wire \u_icache.cblocks[0][31] ;
wire \u_icache.cblocks[0][3] ;
wire \u_icache.cblocks[0][4] ;
wire \u_icache.cblocks[0][5] ;
wire \u_icache.cblocks[0][6] ;
wire \u_icache.cblocks[0][7] ;
wire \u_icache.cblocks[0][8] ;
wire \u_icache.cblocks[0][9] ;
wire \u_icache.cblocks[1][0] ;
wire \u_icache.cblocks[1][10] ;
wire \u_icache.cblocks[1][11] ;
wire \u_icache.cblocks[1][12] ;
wire \u_icache.cblocks[1][13] ;
wire \u_icache.cblocks[1][14] ;
wire \u_icache.cblocks[1][15] ;
wire \u_icache.cblocks[1][16] ;
wire \u_icache.cblocks[1][17] ;
wire \u_icache.cblocks[1][18] ;
wire \u_icache.cblocks[1][19] ;
wire \u_icache.cblocks[1][1] ;
wire \u_icache.cblocks[1][20] ;
wire \u_icache.cblocks[1][21] ;
wire \u_icache.cblocks[1][22] ;
wire \u_icache.cblocks[1][23] ;
wire \u_icache.cblocks[1][24] ;
wire \u_icache.cblocks[1][25] ;
wire \u_icache.cblocks[1][26] ;
wire \u_icache.cblocks[1][27] ;
wire \u_icache.cblocks[1][28] ;
wire \u_icache.cblocks[1][29] ;
wire \u_icache.cblocks[1][2] ;
wire \u_icache.cblocks[1][30] ;
wire \u_icache.cblocks[1][31] ;
wire \u_icache.cblocks[1][3] ;
wire \u_icache.cblocks[1][4] ;
wire \u_icache.cblocks[1][5] ;
wire \u_icache.cblocks[1][6] ;
wire \u_icache.cblocks[1][7] ;
wire \u_icache.cblocks[1][8] ;
wire \u_icache.cblocks[1][9] ;
wire \u_icache.cblocks[2][0] ;
wire \u_icache.cblocks[2][10] ;
wire \u_icache.cblocks[2][11] ;
wire \u_icache.cblocks[2][12] ;
wire \u_icache.cblocks[2][13] ;
wire \u_icache.cblocks[2][14] ;
wire \u_icache.cblocks[2][15] ;
wire \u_icache.cblocks[2][16] ;
wire \u_icache.cblocks[2][17] ;
wire \u_icache.cblocks[2][18] ;
wire \u_icache.cblocks[2][19] ;
wire \u_icache.cblocks[2][1] ;
wire \u_icache.cblocks[2][20] ;
wire \u_icache.cblocks[2][21] ;
wire \u_icache.cblocks[2][22] ;
wire \u_icache.cblocks[2][23] ;
wire \u_icache.cblocks[2][24] ;
wire \u_icache.cblocks[2][25] ;
wire \u_icache.cblocks[2][26] ;
wire \u_icache.cblocks[2][27] ;
wire \u_icache.cblocks[2][28] ;
wire \u_icache.cblocks[2][29] ;
wire \u_icache.cblocks[2][2] ;
wire \u_icache.cblocks[2][30] ;
wire \u_icache.cblocks[2][31] ;
wire \u_icache.cblocks[2][3] ;
wire \u_icache.cblocks[2][4] ;
wire \u_icache.cblocks[2][5] ;
wire \u_icache.cblocks[2][6] ;
wire \u_icache.cblocks[2][7] ;
wire \u_icache.cblocks[2][8] ;
wire \u_icache.cblocks[2][9] ;
wire \u_icache.cblocks[3][0] ;
wire \u_icache.cblocks[3][10] ;
wire \u_icache.cblocks[3][11] ;
wire \u_icache.cblocks[3][12] ;
wire \u_icache.cblocks[3][13] ;
wire \u_icache.cblocks[3][14] ;
wire \u_icache.cblocks[3][15] ;
wire \u_icache.cblocks[3][16] ;
wire \u_icache.cblocks[3][17] ;
wire \u_icache.cblocks[3][18] ;
wire \u_icache.cblocks[3][19] ;
wire \u_icache.cblocks[3][1] ;
wire \u_icache.cblocks[3][20] ;
wire \u_icache.cblocks[3][21] ;
wire \u_icache.cblocks[3][22] ;
wire \u_icache.cblocks[3][23] ;
wire \u_icache.cblocks[3][24] ;
wire \u_icache.cblocks[3][25] ;
wire \u_icache.cblocks[3][26] ;
wire \u_icache.cblocks[3][27] ;
wire \u_icache.cblocks[3][28] ;
wire \u_icache.cblocks[3][29] ;
wire \u_icache.cblocks[3][2] ;
wire \u_icache.cblocks[3][30] ;
wire \u_icache.cblocks[3][31] ;
wire \u_icache.cblocks[3][3] ;
wire \u_icache.cblocks[3][4] ;
wire \u_icache.cblocks[3][5] ;
wire \u_icache.cblocks[3][6] ;
wire \u_icache.cblocks[3][7] ;
wire \u_icache.cblocks[3][8] ;
wire \u_icache.cblocks[3][9] ;
wire \u_icache.cblocks[4][0] ;
wire \u_icache.cblocks[4][10] ;
wire \u_icache.cblocks[4][11] ;
wire \u_icache.cblocks[4][12] ;
wire \u_icache.cblocks[4][13] ;
wire \u_icache.cblocks[4][14] ;
wire \u_icache.cblocks[4][15] ;
wire \u_icache.cblocks[4][16] ;
wire \u_icache.cblocks[4][17] ;
wire \u_icache.cblocks[4][18] ;
wire \u_icache.cblocks[4][19] ;
wire \u_icache.cblocks[4][1] ;
wire \u_icache.cblocks[4][20] ;
wire \u_icache.cblocks[4][21] ;
wire \u_icache.cblocks[4][22] ;
wire \u_icache.cblocks[4][23] ;
wire \u_icache.cblocks[4][24] ;
wire \u_icache.cblocks[4][25] ;
wire \u_icache.cblocks[4][26] ;
wire \u_icache.cblocks[4][27] ;
wire \u_icache.cblocks[4][28] ;
wire \u_icache.cblocks[4][29] ;
wire \u_icache.cblocks[4][2] ;
wire \u_icache.cblocks[4][30] ;
wire \u_icache.cblocks[4][31] ;
wire \u_icache.cblocks[4][3] ;
wire \u_icache.cblocks[4][4] ;
wire \u_icache.cblocks[4][5] ;
wire \u_icache.cblocks[4][6] ;
wire \u_icache.cblocks[4][7] ;
wire \u_icache.cblocks[4][8] ;
wire \u_icache.cblocks[4][9] ;
wire \u_icache.cblocks[5][0] ;
wire \u_icache.cblocks[5][10] ;
wire \u_icache.cblocks[5][11] ;
wire \u_icache.cblocks[5][12] ;
wire \u_icache.cblocks[5][13] ;
wire \u_icache.cblocks[5][14] ;
wire \u_icache.cblocks[5][15] ;
wire \u_icache.cblocks[5][16] ;
wire \u_icache.cblocks[5][17] ;
wire \u_icache.cblocks[5][18] ;
wire \u_icache.cblocks[5][19] ;
wire \u_icache.cblocks[5][1] ;
wire \u_icache.cblocks[5][20] ;
wire \u_icache.cblocks[5][21] ;
wire \u_icache.cblocks[5][22] ;
wire \u_icache.cblocks[5][23] ;
wire \u_icache.cblocks[5][24] ;
wire \u_icache.cblocks[5][25] ;
wire \u_icache.cblocks[5][26] ;
wire \u_icache.cblocks[5][27] ;
wire \u_icache.cblocks[5][28] ;
wire \u_icache.cblocks[5][29] ;
wire \u_icache.cblocks[5][2] ;
wire \u_icache.cblocks[5][30] ;
wire \u_icache.cblocks[5][31] ;
wire \u_icache.cblocks[5][3] ;
wire \u_icache.cblocks[5][4] ;
wire \u_icache.cblocks[5][5] ;
wire \u_icache.cblocks[5][6] ;
wire \u_icache.cblocks[5][7] ;
wire \u_icache.cblocks[5][8] ;
wire \u_icache.cblocks[5][9] ;
wire \u_icache.cblocks[6][0] ;
wire \u_icache.cblocks[6][10] ;
wire \u_icache.cblocks[6][11] ;
wire \u_icache.cblocks[6][12] ;
wire \u_icache.cblocks[6][13] ;
wire \u_icache.cblocks[6][14] ;
wire \u_icache.cblocks[6][15] ;
wire \u_icache.cblocks[6][16] ;
wire \u_icache.cblocks[6][17] ;
wire \u_icache.cblocks[6][18] ;
wire \u_icache.cblocks[6][19] ;
wire \u_icache.cblocks[6][1] ;
wire \u_icache.cblocks[6][20] ;
wire \u_icache.cblocks[6][21] ;
wire \u_icache.cblocks[6][22] ;
wire \u_icache.cblocks[6][23] ;
wire \u_icache.cblocks[6][24] ;
wire \u_icache.cblocks[6][25] ;
wire \u_icache.cblocks[6][26] ;
wire \u_icache.cblocks[6][27] ;
wire \u_icache.cblocks[6][28] ;
wire \u_icache.cblocks[6][29] ;
wire \u_icache.cblocks[6][2] ;
wire \u_icache.cblocks[6][30] ;
wire \u_icache.cblocks[6][31] ;
wire \u_icache.cblocks[6][3] ;
wire \u_icache.cblocks[6][4] ;
wire \u_icache.cblocks[6][5] ;
wire \u_icache.cblocks[6][6] ;
wire \u_icache.cblocks[6][7] ;
wire \u_icache.cblocks[6][8] ;
wire \u_icache.cblocks[6][9] ;
wire \u_icache.cblocks[7][0] ;
wire \u_icache.cblocks[7][10] ;
wire \u_icache.cblocks[7][11] ;
wire \u_icache.cblocks[7][12] ;
wire \u_icache.cblocks[7][13] ;
wire \u_icache.cblocks[7][14] ;
wire \u_icache.cblocks[7][15] ;
wire \u_icache.cblocks[7][16] ;
wire \u_icache.cblocks[7][17] ;
wire \u_icache.cblocks[7][18] ;
wire \u_icache.cblocks[7][19] ;
wire \u_icache.cblocks[7][1] ;
wire \u_icache.cblocks[7][20] ;
wire \u_icache.cblocks[7][21] ;
wire \u_icache.cblocks[7][22] ;
wire \u_icache.cblocks[7][23] ;
wire \u_icache.cblocks[7][24] ;
wire \u_icache.cblocks[7][25] ;
wire \u_icache.cblocks[7][26] ;
wire \u_icache.cblocks[7][27] ;
wire \u_icache.cblocks[7][28] ;
wire \u_icache.cblocks[7][29] ;
wire \u_icache.cblocks[7][2] ;
wire \u_icache.cblocks[7][30] ;
wire \u_icache.cblocks[7][31] ;
wire \u_icache.cblocks[7][3] ;
wire \u_icache.cblocks[7][4] ;
wire \u_icache.cblocks[7][5] ;
wire \u_icache.cblocks[7][6] ;
wire \u_icache.cblocks[7][7] ;
wire \u_icache.cblocks[7][8] ;
wire \u_icache.cblocks[7][9] ;
wire \u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ;
wire \u_icache.chvalid_$_SDFFE_PP0P__Q_E ;
wire \u_icache.count_$_NOT__A_Y ;
wire \u_icache.count_$_SDFFE_PP0P__Q_E ;
wire \u_icache.cready_$_ANDNOT__A_Y ;
wire \u_icache.cready_$_ANDNOT__B_Y_$_OR__B_Y ;
wire \u_icache.ctags[0][0] ;
wire \u_icache.ctags[0][10] ;
wire \u_icache.ctags[0][11] ;
wire \u_icache.ctags[0][12] ;
wire \u_icache.ctags[0][13] ;
wire \u_icache.ctags[0][14] ;
wire \u_icache.ctags[0][15] ;
wire \u_icache.ctags[0][16] ;
wire \u_icache.ctags[0][17] ;
wire \u_icache.ctags[0][18] ;
wire \u_icache.ctags[0][19] ;
wire \u_icache.ctags[0][1] ;
wire \u_icache.ctags[0][20] ;
wire \u_icache.ctags[0][21] ;
wire \u_icache.ctags[0][22] ;
wire \u_icache.ctags[0][23] ;
wire \u_icache.ctags[0][24] ;
wire \u_icache.ctags[0][25] ;
wire \u_icache.ctags[0][26] ;
wire \u_icache.ctags[0][2] ;
wire \u_icache.ctags[0][3] ;
wire \u_icache.ctags[0][4] ;
wire \u_icache.ctags[0][5] ;
wire \u_icache.ctags[0][6] ;
wire \u_icache.ctags[0][7] ;
wire \u_icache.ctags[0][8] ;
wire \u_icache.ctags[0][9] ;
wire \u_icache.ctags[1][0] ;
wire \u_icache.ctags[1][10] ;
wire \u_icache.ctags[1][11] ;
wire \u_icache.ctags[1][12] ;
wire \u_icache.ctags[1][13] ;
wire \u_icache.ctags[1][14] ;
wire \u_icache.ctags[1][15] ;
wire \u_icache.ctags[1][16] ;
wire \u_icache.ctags[1][17] ;
wire \u_icache.ctags[1][18] ;
wire \u_icache.ctags[1][19] ;
wire \u_icache.ctags[1][1] ;
wire \u_icache.ctags[1][20] ;
wire \u_icache.ctags[1][21] ;
wire \u_icache.ctags[1][22] ;
wire \u_icache.ctags[1][23] ;
wire \u_icache.ctags[1][24] ;
wire \u_icache.ctags[1][25] ;
wire \u_icache.ctags[1][26] ;
wire \u_icache.ctags[1][2] ;
wire \u_icache.ctags[1][3] ;
wire \u_icache.ctags[1][4] ;
wire \u_icache.ctags[1][5] ;
wire \u_icache.ctags[1][6] ;
wire \u_icache.ctags[1][7] ;
wire \u_icache.ctags[1][8] ;
wire \u_icache.ctags[1][9] ;
wire \u_icache.cvalids_$_SDFFE_PP0P__Q_E ;
wire \u_icache.ended ;
wire \u_icache.ended_$_ANDNOT__B_Y ;
wire \u_icache.ended_$_SDFFE_PP0P__Q_E ;
wire \u_idu.decode_ok_$_SDFFE_PP0P__Q_E ;
wire \u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ;
wire \u_ifu.inst_ok_$_ANDNOT__A_Y ;
wire \u_ifu.inst_ok_$_SDFFE_PP0P__Q_E ;
wire \u_ifu.jpc_ok ;
wire \u_ifu.jpc_ok_$_NOT__A_Y ;
wire \u_ifu.jpc_ok_$_SDFFE_PP0P__Q_E ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_B_$_ANDNOT__B_Y ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_Y ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_28_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_ifu.pc_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.arvalid ;
wire \u_lsu.arvalid_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.awvalid_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.reading ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_1_Y ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_2_Y ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_3_Y ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_4_Y ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_5_Y ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_6_Y ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_7_Y ;
wire \u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ;
wire \u_lsu.reading_$_NOR__B_A_$_MUX__Y_A ;
wire \u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ;
wire \u_lsu.reading_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.rvalid ;
wire \u_lsu.rvalid_clint ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_10_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_18_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_26_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_28_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_31_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_39_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_8_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ;
wire \u_lsu.wlast_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.writing ;
wire \u_reg.rf[10][0] ;
wire \u_reg.rf[10][10] ;
wire \u_reg.rf[10][11] ;
wire \u_reg.rf[10][12] ;
wire \u_reg.rf[10][13] ;
wire \u_reg.rf[10][14] ;
wire \u_reg.rf[10][15] ;
wire \u_reg.rf[10][16] ;
wire \u_reg.rf[10][17] ;
wire \u_reg.rf[10][18] ;
wire \u_reg.rf[10][19] ;
wire \u_reg.rf[10][1] ;
wire \u_reg.rf[10][20] ;
wire \u_reg.rf[10][21] ;
wire \u_reg.rf[10][22] ;
wire \u_reg.rf[10][23] ;
wire \u_reg.rf[10][24] ;
wire \u_reg.rf[10][25] ;
wire \u_reg.rf[10][26] ;
wire \u_reg.rf[10][27] ;
wire \u_reg.rf[10][28] ;
wire \u_reg.rf[10][29] ;
wire \u_reg.rf[10][2] ;
wire \u_reg.rf[10][30] ;
wire \u_reg.rf[10][31] ;
wire \u_reg.rf[10][3] ;
wire \u_reg.rf[10][4] ;
wire \u_reg.rf[10][5] ;
wire \u_reg.rf[10][6] ;
wire \u_reg.rf[10][7] ;
wire \u_reg.rf[10][8] ;
wire \u_reg.rf[10][9] ;
wire \u_reg.rf[11][0] ;
wire \u_reg.rf[11][10] ;
wire \u_reg.rf[11][11] ;
wire \u_reg.rf[11][12] ;
wire \u_reg.rf[11][13] ;
wire \u_reg.rf[11][14] ;
wire \u_reg.rf[11][15] ;
wire \u_reg.rf[11][16] ;
wire \u_reg.rf[11][17] ;
wire \u_reg.rf[11][18] ;
wire \u_reg.rf[11][19] ;
wire \u_reg.rf[11][1] ;
wire \u_reg.rf[11][20] ;
wire \u_reg.rf[11][21] ;
wire \u_reg.rf[11][22] ;
wire \u_reg.rf[11][23] ;
wire \u_reg.rf[11][24] ;
wire \u_reg.rf[11][25] ;
wire \u_reg.rf[11][26] ;
wire \u_reg.rf[11][27] ;
wire \u_reg.rf[11][28] ;
wire \u_reg.rf[11][29] ;
wire \u_reg.rf[11][2] ;
wire \u_reg.rf[11][30] ;
wire \u_reg.rf[11][31] ;
wire \u_reg.rf[11][3] ;
wire \u_reg.rf[11][4] ;
wire \u_reg.rf[11][5] ;
wire \u_reg.rf[11][6] ;
wire \u_reg.rf[11][7] ;
wire \u_reg.rf[11][8] ;
wire \u_reg.rf[11][9] ;
wire \u_reg.rf[12][0] ;
wire \u_reg.rf[12][10] ;
wire \u_reg.rf[12][11] ;
wire \u_reg.rf[12][12] ;
wire \u_reg.rf[12][13] ;
wire \u_reg.rf[12][14] ;
wire \u_reg.rf[12][15] ;
wire \u_reg.rf[12][16] ;
wire \u_reg.rf[12][17] ;
wire \u_reg.rf[12][18] ;
wire \u_reg.rf[12][19] ;
wire \u_reg.rf[12][1] ;
wire \u_reg.rf[12][20] ;
wire \u_reg.rf[12][21] ;
wire \u_reg.rf[12][22] ;
wire \u_reg.rf[12][23] ;
wire \u_reg.rf[12][24] ;
wire \u_reg.rf[12][25] ;
wire \u_reg.rf[12][26] ;
wire \u_reg.rf[12][27] ;
wire \u_reg.rf[12][28] ;
wire \u_reg.rf[12][29] ;
wire \u_reg.rf[12][2] ;
wire \u_reg.rf[12][30] ;
wire \u_reg.rf[12][31] ;
wire \u_reg.rf[12][3] ;
wire \u_reg.rf[12][4] ;
wire \u_reg.rf[12][5] ;
wire \u_reg.rf[12][6] ;
wire \u_reg.rf[12][7] ;
wire \u_reg.rf[12][8] ;
wire \u_reg.rf[12][9] ;
wire \u_reg.rf[13][0] ;
wire \u_reg.rf[13][10] ;
wire \u_reg.rf[13][11] ;
wire \u_reg.rf[13][12] ;
wire \u_reg.rf[13][13] ;
wire \u_reg.rf[13][14] ;
wire \u_reg.rf[13][15] ;
wire \u_reg.rf[13][16] ;
wire \u_reg.rf[13][17] ;
wire \u_reg.rf[13][18] ;
wire \u_reg.rf[13][19] ;
wire \u_reg.rf[13][1] ;
wire \u_reg.rf[13][20] ;
wire \u_reg.rf[13][21] ;
wire \u_reg.rf[13][22] ;
wire \u_reg.rf[13][23] ;
wire \u_reg.rf[13][24] ;
wire \u_reg.rf[13][25] ;
wire \u_reg.rf[13][26] ;
wire \u_reg.rf[13][27] ;
wire \u_reg.rf[13][28] ;
wire \u_reg.rf[13][29] ;
wire \u_reg.rf[13][2] ;
wire \u_reg.rf[13][30] ;
wire \u_reg.rf[13][31] ;
wire \u_reg.rf[13][3] ;
wire \u_reg.rf[13][4] ;
wire \u_reg.rf[13][5] ;
wire \u_reg.rf[13][6] ;
wire \u_reg.rf[13][7] ;
wire \u_reg.rf[13][8] ;
wire \u_reg.rf[13][9] ;
wire \u_reg.rf[14][0] ;
wire \u_reg.rf[14][10] ;
wire \u_reg.rf[14][11] ;
wire \u_reg.rf[14][12] ;
wire \u_reg.rf[14][13] ;
wire \u_reg.rf[14][14] ;
wire \u_reg.rf[14][15] ;
wire \u_reg.rf[14][16] ;
wire \u_reg.rf[14][17] ;
wire \u_reg.rf[14][18] ;
wire \u_reg.rf[14][19] ;
wire \u_reg.rf[14][1] ;
wire \u_reg.rf[14][20] ;
wire \u_reg.rf[14][21] ;
wire \u_reg.rf[14][22] ;
wire \u_reg.rf[14][23] ;
wire \u_reg.rf[14][24] ;
wire \u_reg.rf[14][25] ;
wire \u_reg.rf[14][26] ;
wire \u_reg.rf[14][27] ;
wire \u_reg.rf[14][28] ;
wire \u_reg.rf[14][29] ;
wire \u_reg.rf[14][2] ;
wire \u_reg.rf[14][30] ;
wire \u_reg.rf[14][31] ;
wire \u_reg.rf[14][3] ;
wire \u_reg.rf[14][4] ;
wire \u_reg.rf[14][5] ;
wire \u_reg.rf[14][6] ;
wire \u_reg.rf[14][7] ;
wire \u_reg.rf[14][8] ;
wire \u_reg.rf[14][9] ;
wire \u_reg.rf[15][0] ;
wire \u_reg.rf[15][10] ;
wire \u_reg.rf[15][11] ;
wire \u_reg.rf[15][12] ;
wire \u_reg.rf[15][13] ;
wire \u_reg.rf[15][14] ;
wire \u_reg.rf[15][15] ;
wire \u_reg.rf[15][16] ;
wire \u_reg.rf[15][17] ;
wire \u_reg.rf[15][18] ;
wire \u_reg.rf[15][19] ;
wire \u_reg.rf[15][1] ;
wire \u_reg.rf[15][20] ;
wire \u_reg.rf[15][21] ;
wire \u_reg.rf[15][22] ;
wire \u_reg.rf[15][23] ;
wire \u_reg.rf[15][24] ;
wire \u_reg.rf[15][25] ;
wire \u_reg.rf[15][26] ;
wire \u_reg.rf[15][27] ;
wire \u_reg.rf[15][28] ;
wire \u_reg.rf[15][29] ;
wire \u_reg.rf[15][2] ;
wire \u_reg.rf[15][30] ;
wire \u_reg.rf[15][31] ;
wire \u_reg.rf[15][3] ;
wire \u_reg.rf[15][4] ;
wire \u_reg.rf[15][5] ;
wire \u_reg.rf[15][6] ;
wire \u_reg.rf[15][7] ;
wire \u_reg.rf[15][8] ;
wire \u_reg.rf[15][9] ;
wire \u_reg.rf[1][0] ;
wire \u_reg.rf[1][10] ;
wire \u_reg.rf[1][11] ;
wire \u_reg.rf[1][12] ;
wire \u_reg.rf[1][13] ;
wire \u_reg.rf[1][14] ;
wire \u_reg.rf[1][15] ;
wire \u_reg.rf[1][16] ;
wire \u_reg.rf[1][17] ;
wire \u_reg.rf[1][18] ;
wire \u_reg.rf[1][19] ;
wire \u_reg.rf[1][1] ;
wire \u_reg.rf[1][20] ;
wire \u_reg.rf[1][21] ;
wire \u_reg.rf[1][22] ;
wire \u_reg.rf[1][23] ;
wire \u_reg.rf[1][24] ;
wire \u_reg.rf[1][25] ;
wire \u_reg.rf[1][26] ;
wire \u_reg.rf[1][27] ;
wire \u_reg.rf[1][28] ;
wire \u_reg.rf[1][29] ;
wire \u_reg.rf[1][2] ;
wire \u_reg.rf[1][30] ;
wire \u_reg.rf[1][31] ;
wire \u_reg.rf[1][3] ;
wire \u_reg.rf[1][4] ;
wire \u_reg.rf[1][5] ;
wire \u_reg.rf[1][6] ;
wire \u_reg.rf[1][7] ;
wire \u_reg.rf[1][8] ;
wire \u_reg.rf[1][9] ;
wire \u_reg.rf[2][0] ;
wire \u_reg.rf[2][10] ;
wire \u_reg.rf[2][11] ;
wire \u_reg.rf[2][12] ;
wire \u_reg.rf[2][13] ;
wire \u_reg.rf[2][14] ;
wire \u_reg.rf[2][15] ;
wire \u_reg.rf[2][16] ;
wire \u_reg.rf[2][17] ;
wire \u_reg.rf[2][18] ;
wire \u_reg.rf[2][19] ;
wire \u_reg.rf[2][1] ;
wire \u_reg.rf[2][20] ;
wire \u_reg.rf[2][21] ;
wire \u_reg.rf[2][22] ;
wire \u_reg.rf[2][23] ;
wire \u_reg.rf[2][24] ;
wire \u_reg.rf[2][25] ;
wire \u_reg.rf[2][26] ;
wire \u_reg.rf[2][27] ;
wire \u_reg.rf[2][28] ;
wire \u_reg.rf[2][29] ;
wire \u_reg.rf[2][2] ;
wire \u_reg.rf[2][30] ;
wire \u_reg.rf[2][31] ;
wire \u_reg.rf[2][3] ;
wire \u_reg.rf[2][4] ;
wire \u_reg.rf[2][5] ;
wire \u_reg.rf[2][6] ;
wire \u_reg.rf[2][7] ;
wire \u_reg.rf[2][8] ;
wire \u_reg.rf[2][9] ;
wire \u_reg.rf[3][0] ;
wire \u_reg.rf[3][10] ;
wire \u_reg.rf[3][11] ;
wire \u_reg.rf[3][12] ;
wire \u_reg.rf[3][13] ;
wire \u_reg.rf[3][14] ;
wire \u_reg.rf[3][15] ;
wire \u_reg.rf[3][16] ;
wire \u_reg.rf[3][17] ;
wire \u_reg.rf[3][18] ;
wire \u_reg.rf[3][19] ;
wire \u_reg.rf[3][1] ;
wire \u_reg.rf[3][20] ;
wire \u_reg.rf[3][21] ;
wire \u_reg.rf[3][22] ;
wire \u_reg.rf[3][23] ;
wire \u_reg.rf[3][24] ;
wire \u_reg.rf[3][25] ;
wire \u_reg.rf[3][26] ;
wire \u_reg.rf[3][27] ;
wire \u_reg.rf[3][28] ;
wire \u_reg.rf[3][29] ;
wire \u_reg.rf[3][2] ;
wire \u_reg.rf[3][30] ;
wire \u_reg.rf[3][31] ;
wire \u_reg.rf[3][3] ;
wire \u_reg.rf[3][4] ;
wire \u_reg.rf[3][5] ;
wire \u_reg.rf[3][6] ;
wire \u_reg.rf[3][7] ;
wire \u_reg.rf[3][8] ;
wire \u_reg.rf[3][9] ;
wire \u_reg.rf[4][0] ;
wire \u_reg.rf[4][10] ;
wire \u_reg.rf[4][11] ;
wire \u_reg.rf[4][12] ;
wire \u_reg.rf[4][13] ;
wire \u_reg.rf[4][14] ;
wire \u_reg.rf[4][15] ;
wire \u_reg.rf[4][16] ;
wire \u_reg.rf[4][17] ;
wire \u_reg.rf[4][18] ;
wire \u_reg.rf[4][19] ;
wire \u_reg.rf[4][1] ;
wire \u_reg.rf[4][20] ;
wire \u_reg.rf[4][21] ;
wire \u_reg.rf[4][22] ;
wire \u_reg.rf[4][23] ;
wire \u_reg.rf[4][24] ;
wire \u_reg.rf[4][25] ;
wire \u_reg.rf[4][26] ;
wire \u_reg.rf[4][27] ;
wire \u_reg.rf[4][28] ;
wire \u_reg.rf[4][29] ;
wire \u_reg.rf[4][2] ;
wire \u_reg.rf[4][30] ;
wire \u_reg.rf[4][31] ;
wire \u_reg.rf[4][3] ;
wire \u_reg.rf[4][4] ;
wire \u_reg.rf[4][5] ;
wire \u_reg.rf[4][6] ;
wire \u_reg.rf[4][7] ;
wire \u_reg.rf[4][8] ;
wire \u_reg.rf[4][9] ;
wire \u_reg.rf[5][0] ;
wire \u_reg.rf[5][10] ;
wire \u_reg.rf[5][11] ;
wire \u_reg.rf[5][12] ;
wire \u_reg.rf[5][13] ;
wire \u_reg.rf[5][14] ;
wire \u_reg.rf[5][15] ;
wire \u_reg.rf[5][16] ;
wire \u_reg.rf[5][17] ;
wire \u_reg.rf[5][18] ;
wire \u_reg.rf[5][19] ;
wire \u_reg.rf[5][1] ;
wire \u_reg.rf[5][20] ;
wire \u_reg.rf[5][21] ;
wire \u_reg.rf[5][22] ;
wire \u_reg.rf[5][23] ;
wire \u_reg.rf[5][24] ;
wire \u_reg.rf[5][25] ;
wire \u_reg.rf[5][26] ;
wire \u_reg.rf[5][27] ;
wire \u_reg.rf[5][28] ;
wire \u_reg.rf[5][29] ;
wire \u_reg.rf[5][2] ;
wire \u_reg.rf[5][30] ;
wire \u_reg.rf[5][31] ;
wire \u_reg.rf[5][3] ;
wire \u_reg.rf[5][4] ;
wire \u_reg.rf[5][5] ;
wire \u_reg.rf[5][6] ;
wire \u_reg.rf[5][7] ;
wire \u_reg.rf[5][8] ;
wire \u_reg.rf[5][9] ;
wire \u_reg.rf[6][0] ;
wire \u_reg.rf[6][10] ;
wire \u_reg.rf[6][11] ;
wire \u_reg.rf[6][12] ;
wire \u_reg.rf[6][13] ;
wire \u_reg.rf[6][14] ;
wire \u_reg.rf[6][15] ;
wire \u_reg.rf[6][16] ;
wire \u_reg.rf[6][17] ;
wire \u_reg.rf[6][18] ;
wire \u_reg.rf[6][19] ;
wire \u_reg.rf[6][1] ;
wire \u_reg.rf[6][20] ;
wire \u_reg.rf[6][21] ;
wire \u_reg.rf[6][22] ;
wire \u_reg.rf[6][23] ;
wire \u_reg.rf[6][24] ;
wire \u_reg.rf[6][25] ;
wire \u_reg.rf[6][26] ;
wire \u_reg.rf[6][27] ;
wire \u_reg.rf[6][28] ;
wire \u_reg.rf[6][29] ;
wire \u_reg.rf[6][2] ;
wire \u_reg.rf[6][30] ;
wire \u_reg.rf[6][31] ;
wire \u_reg.rf[6][3] ;
wire \u_reg.rf[6][4] ;
wire \u_reg.rf[6][5] ;
wire \u_reg.rf[6][6] ;
wire \u_reg.rf[6][7] ;
wire \u_reg.rf[6][8] ;
wire \u_reg.rf[6][9] ;
wire \u_reg.rf[7][0] ;
wire \u_reg.rf[7][10] ;
wire \u_reg.rf[7][11] ;
wire \u_reg.rf[7][12] ;
wire \u_reg.rf[7][13] ;
wire \u_reg.rf[7][14] ;
wire \u_reg.rf[7][15] ;
wire \u_reg.rf[7][16] ;
wire \u_reg.rf[7][17] ;
wire \u_reg.rf[7][18] ;
wire \u_reg.rf[7][19] ;
wire \u_reg.rf[7][1] ;
wire \u_reg.rf[7][20] ;
wire \u_reg.rf[7][21] ;
wire \u_reg.rf[7][22] ;
wire \u_reg.rf[7][23] ;
wire \u_reg.rf[7][24] ;
wire \u_reg.rf[7][25] ;
wire \u_reg.rf[7][26] ;
wire \u_reg.rf[7][27] ;
wire \u_reg.rf[7][28] ;
wire \u_reg.rf[7][29] ;
wire \u_reg.rf[7][2] ;
wire \u_reg.rf[7][30] ;
wire \u_reg.rf[7][31] ;
wire \u_reg.rf[7][3] ;
wire \u_reg.rf[7][4] ;
wire \u_reg.rf[7][5] ;
wire \u_reg.rf[7][6] ;
wire \u_reg.rf[7][7] ;
wire \u_reg.rf[7][8] ;
wire \u_reg.rf[7][9] ;
wire \u_reg.rf[8][0] ;
wire \u_reg.rf[8][10] ;
wire \u_reg.rf[8][11] ;
wire \u_reg.rf[8][12] ;
wire \u_reg.rf[8][13] ;
wire \u_reg.rf[8][14] ;
wire \u_reg.rf[8][15] ;
wire \u_reg.rf[8][16] ;
wire \u_reg.rf[8][17] ;
wire \u_reg.rf[8][18] ;
wire \u_reg.rf[8][19] ;
wire \u_reg.rf[8][1] ;
wire \u_reg.rf[8][20] ;
wire \u_reg.rf[8][21] ;
wire \u_reg.rf[8][22] ;
wire \u_reg.rf[8][23] ;
wire \u_reg.rf[8][24] ;
wire \u_reg.rf[8][25] ;
wire \u_reg.rf[8][26] ;
wire \u_reg.rf[8][27] ;
wire \u_reg.rf[8][28] ;
wire \u_reg.rf[8][29] ;
wire \u_reg.rf[8][2] ;
wire \u_reg.rf[8][30] ;
wire \u_reg.rf[8][31] ;
wire \u_reg.rf[8][3] ;
wire \u_reg.rf[8][4] ;
wire \u_reg.rf[8][5] ;
wire \u_reg.rf[8][6] ;
wire \u_reg.rf[8][7] ;
wire \u_reg.rf[8][8] ;
wire \u_reg.rf[8][9] ;
wire \u_reg.rf[9][0] ;
wire \u_reg.rf[9][10] ;
wire \u_reg.rf[9][11] ;
wire \u_reg.rf[9][12] ;
wire \u_reg.rf[9][13] ;
wire \u_reg.rf[9][14] ;
wire \u_reg.rf[9][15] ;
wire \u_reg.rf[9][16] ;
wire \u_reg.rf[9][17] ;
wire \u_reg.rf[9][18] ;
wire \u_reg.rf[9][19] ;
wire \u_reg.rf[9][1] ;
wire \u_reg.rf[9][20] ;
wire \u_reg.rf[9][21] ;
wire \u_reg.rf[9][22] ;
wire \u_reg.rf[9][23] ;
wire \u_reg.rf[9][24] ;
wire \u_reg.rf[9][25] ;
wire \u_reg.rf[9][26] ;
wire \u_reg.rf[9][27] ;
wire \u_reg.rf[9][28] ;
wire \u_reg.rf[9][29] ;
wire \u_reg.rf[9][2] ;
wire \u_reg.rf[9][30] ;
wire \u_reg.rf[9][31] ;
wire \u_reg.rf[9][3] ;
wire \u_reg.rf[9][4] ;
wire \u_reg.rf[9][5] ;
wire \u_reg.rf[9][6] ;
wire \u_reg.rf[9][7] ;
wire \u_reg.rf[9][8] ;
wire \u_reg.rf[9][9] ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire \io_master_awaddr[0] ;
wire \io_master_awaddr[1] ;
wire \io_master_awaddr[2] ;
wire \io_master_awaddr[3] ;
wire \io_master_awaddr[4] ;
wire \io_master_awaddr[5] ;
wire \io_master_awaddr[6] ;
wire \io_master_awaddr[7] ;
wire \io_master_awaddr[8] ;
wire \io_master_awaddr[9] ;
wire \io_master_awaddr[10] ;
wire \io_master_awaddr[11] ;
wire \io_master_awaddr[12] ;
wire \io_master_awaddr[13] ;
wire \io_master_awaddr[14] ;
wire \io_master_awaddr[15] ;
wire \io_master_awaddr[16] ;
wire \io_master_awaddr[17] ;
wire \io_master_awaddr[18] ;
wire \io_master_awaddr[19] ;
wire \io_master_awaddr[20] ;
wire \io_master_awaddr[21] ;
wire \io_master_awaddr[22] ;
wire \io_master_awaddr[23] ;
wire \io_master_awaddr[24] ;
wire \io_master_awaddr[25] ;
wire \io_master_awaddr[26] ;
wire \io_master_awaddr[27] ;
wire \io_master_awaddr[28] ;
wire \io_master_awaddr[29] ;
wire \io_master_awaddr[30] ;
wire \io_master_awaddr[31] ;
wire \io_master_awid[0] ;
wire \io_master_awid[1] ;
wire \io_master_awid[2] ;
wire \io_master_awid[3] ;
wire \io_master_awlen[0] ;
wire \io_master_awlen[1] ;
wire \io_master_awlen[2] ;
wire \io_master_awlen[3] ;
wire \io_master_awlen[4] ;
wire \io_master_awlen[5] ;
wire \io_master_awlen[6] ;
wire \io_master_awlen[7] ;
wire \io_master_awsize[0] ;
wire \io_master_awsize[1] ;
wire \io_master_awsize[2] ;
wire \io_master_awburst[0] ;
wire \io_master_awburst[1] ;
wire \io_master_wdata[0] ;
wire \io_master_wdata[1] ;
wire \io_master_wdata[2] ;
wire \io_master_wdata[3] ;
wire \io_master_wdata[4] ;
wire \io_master_wdata[5] ;
wire \io_master_wdata[6] ;
wire \io_master_wdata[7] ;
wire \io_master_wdata[8] ;
wire \io_master_wdata[9] ;
wire \io_master_wdata[10] ;
wire \io_master_wdata[11] ;
wire \io_master_wdata[12] ;
wire \io_master_wdata[13] ;
wire \io_master_wdata[14] ;
wire \io_master_wdata[15] ;
wire \io_master_wdata[16] ;
wire \io_master_wdata[17] ;
wire \io_master_wdata[18] ;
wire \io_master_wdata[19] ;
wire \io_master_wdata[20] ;
wire \io_master_wdata[21] ;
wire \io_master_wdata[22] ;
wire \io_master_wdata[23] ;
wire \io_master_wdata[24] ;
wire \io_master_wdata[25] ;
wire \io_master_wdata[26] ;
wire \io_master_wdata[27] ;
wire \io_master_wdata[28] ;
wire \io_master_wdata[29] ;
wire \io_master_wdata[30] ;
wire \io_master_wdata[31] ;
wire \io_master_wstrb[0] ;
wire \io_master_wstrb[1] ;
wire \io_master_wstrb[2] ;
wire \io_master_wstrb[3] ;
wire \io_master_bresp[0] ;
wire \io_master_bresp[1] ;
wire \io_master_bid[0] ;
wire \io_master_bid[1] ;
wire \io_master_bid[2] ;
wire \io_master_bid[3] ;
wire \io_master_araddr[0] ;
wire \io_master_araddr[1] ;
wire \io_master_araddr[2] ;
wire \io_master_araddr[3] ;
wire \io_master_araddr[4] ;
wire \io_master_araddr[5] ;
wire \io_master_araddr[6] ;
wire \io_master_araddr[7] ;
wire \io_master_araddr[8] ;
wire \io_master_araddr[9] ;
wire \io_master_araddr[10] ;
wire \io_master_araddr[11] ;
wire \io_master_araddr[12] ;
wire \io_master_araddr[13] ;
wire \io_master_araddr[14] ;
wire \io_master_araddr[15] ;
wire \io_master_araddr[16] ;
wire \io_master_araddr[17] ;
wire \io_master_araddr[18] ;
wire \io_master_araddr[19] ;
wire \io_master_araddr[20] ;
wire \io_master_araddr[21] ;
wire \io_master_araddr[22] ;
wire \io_master_araddr[23] ;
wire \io_master_araddr[24] ;
wire \io_master_araddr[25] ;
wire \io_master_araddr[26] ;
wire \io_master_araddr[27] ;
wire \io_master_araddr[28] ;
wire \io_master_araddr[29] ;
wire \io_master_araddr[30] ;
wire \io_master_araddr[31] ;
wire \io_master_arid[0] ;
wire \io_master_arid[1] ;
wire \io_master_arid[2] ;
wire \io_master_arid[3] ;
wire \io_master_arlen[0] ;
wire \io_master_arlen[1] ;
wire \io_master_arlen[2] ;
wire \io_master_arlen[3] ;
wire \io_master_arlen[4] ;
wire \io_master_arlen[5] ;
wire \io_master_arlen[6] ;
wire \io_master_arlen[7] ;
wire \io_master_arsize[0] ;
wire \io_master_arsize[1] ;
wire \io_master_arsize[2] ;
wire \io_master_arburst[0] ;
wire \io_master_arburst[1] ;
wire \io_master_rresp[0] ;
wire \io_master_rresp[1] ;
wire \io_master_rdata[0] ;
wire \io_master_rdata[1] ;
wire \io_master_rdata[2] ;
wire \io_master_rdata[3] ;
wire \io_master_rdata[4] ;
wire \io_master_rdata[5] ;
wire \io_master_rdata[6] ;
wire \io_master_rdata[7] ;
wire \io_master_rdata[8] ;
wire \io_master_rdata[9] ;
wire \io_master_rdata[10] ;
wire \io_master_rdata[11] ;
wire \io_master_rdata[12] ;
wire \io_master_rdata[13] ;
wire \io_master_rdata[14] ;
wire \io_master_rdata[15] ;
wire \io_master_rdata[16] ;
wire \io_master_rdata[17] ;
wire \io_master_rdata[18] ;
wire \io_master_rdata[19] ;
wire \io_master_rdata[20] ;
wire \io_master_rdata[21] ;
wire \io_master_rdata[22] ;
wire \io_master_rdata[23] ;
wire \io_master_rdata[24] ;
wire \io_master_rdata[25] ;
wire \io_master_rdata[26] ;
wire \io_master_rdata[27] ;
wire \io_master_rdata[28] ;
wire \io_master_rdata[29] ;
wire \io_master_rdata[30] ;
wire \io_master_rdata[31] ;
wire \io_master_rid[0] ;
wire \io_master_rid[1] ;
wire \io_master_rid[2] ;
wire \io_master_rid[3] ;
wire \io_slave_awaddr[0] ;
wire \io_slave_awaddr[1] ;
wire \io_slave_awaddr[2] ;
wire \io_slave_awaddr[3] ;
wire \io_slave_awaddr[4] ;
wire \io_slave_awaddr[5] ;
wire \io_slave_awaddr[6] ;
wire \io_slave_awaddr[7] ;
wire \io_slave_awaddr[8] ;
wire \io_slave_awaddr[9] ;
wire \io_slave_awaddr[10] ;
wire \io_slave_awaddr[11] ;
wire \io_slave_awaddr[12] ;
wire \io_slave_awaddr[13] ;
wire \io_slave_awaddr[14] ;
wire \io_slave_awaddr[15] ;
wire \io_slave_awaddr[16] ;
wire \io_slave_awaddr[17] ;
wire \io_slave_awaddr[18] ;
wire \io_slave_awaddr[19] ;
wire \io_slave_awaddr[20] ;
wire \io_slave_awaddr[21] ;
wire \io_slave_awaddr[22] ;
wire \io_slave_awaddr[23] ;
wire \io_slave_awaddr[24] ;
wire \io_slave_awaddr[25] ;
wire \io_slave_awaddr[26] ;
wire \io_slave_awaddr[27] ;
wire \io_slave_awaddr[28] ;
wire \io_slave_awaddr[29] ;
wire \io_slave_awaddr[30] ;
wire \io_slave_awaddr[31] ;
wire \io_slave_awid[0] ;
wire \io_slave_awid[1] ;
wire \io_slave_awid[2] ;
wire \io_slave_awid[3] ;
wire \io_slave_awlen[0] ;
wire \io_slave_awlen[1] ;
wire \io_slave_awlen[2] ;
wire \io_slave_awlen[3] ;
wire \io_slave_awlen[4] ;
wire \io_slave_awlen[5] ;
wire \io_slave_awlen[6] ;
wire \io_slave_awlen[7] ;
wire \io_slave_awsize[0] ;
wire \io_slave_awsize[1] ;
wire \io_slave_awsize[2] ;
wire \io_slave_awburst[0] ;
wire \io_slave_awburst[1] ;
wire \io_slave_wdata[0] ;
wire \io_slave_wdata[1] ;
wire \io_slave_wdata[2] ;
wire \io_slave_wdata[3] ;
wire \io_slave_wdata[4] ;
wire \io_slave_wdata[5] ;
wire \io_slave_wdata[6] ;
wire \io_slave_wdata[7] ;
wire \io_slave_wdata[8] ;
wire \io_slave_wdata[9] ;
wire \io_slave_wdata[10] ;
wire \io_slave_wdata[11] ;
wire \io_slave_wdata[12] ;
wire \io_slave_wdata[13] ;
wire \io_slave_wdata[14] ;
wire \io_slave_wdata[15] ;
wire \io_slave_wdata[16] ;
wire \io_slave_wdata[17] ;
wire \io_slave_wdata[18] ;
wire \io_slave_wdata[19] ;
wire \io_slave_wdata[20] ;
wire \io_slave_wdata[21] ;
wire \io_slave_wdata[22] ;
wire \io_slave_wdata[23] ;
wire \io_slave_wdata[24] ;
wire \io_slave_wdata[25] ;
wire \io_slave_wdata[26] ;
wire \io_slave_wdata[27] ;
wire \io_slave_wdata[28] ;
wire \io_slave_wdata[29] ;
wire \io_slave_wdata[30] ;
wire \io_slave_wdata[31] ;
wire \io_slave_wstrb[0] ;
wire \io_slave_wstrb[1] ;
wire \io_slave_wstrb[2] ;
wire \io_slave_wstrb[3] ;
wire \io_slave_bresp[0] ;
wire \io_slave_bresp[1] ;
wire \io_slave_bid[0] ;
wire \io_slave_bid[1] ;
wire \io_slave_bid[2] ;
wire \io_slave_bid[3] ;
wire \io_slave_araddr[0] ;
wire \io_slave_araddr[1] ;
wire \io_slave_araddr[2] ;
wire \io_slave_araddr[3] ;
wire \io_slave_araddr[4] ;
wire \io_slave_araddr[5] ;
wire \io_slave_araddr[6] ;
wire \io_slave_araddr[7] ;
wire \io_slave_araddr[8] ;
wire \io_slave_araddr[9] ;
wire \io_slave_araddr[10] ;
wire \io_slave_araddr[11] ;
wire \io_slave_araddr[12] ;
wire \io_slave_araddr[13] ;
wire \io_slave_araddr[14] ;
wire \io_slave_araddr[15] ;
wire \io_slave_araddr[16] ;
wire \io_slave_araddr[17] ;
wire \io_slave_araddr[18] ;
wire \io_slave_araddr[19] ;
wire \io_slave_araddr[20] ;
wire \io_slave_araddr[21] ;
wire \io_slave_araddr[22] ;
wire \io_slave_araddr[23] ;
wire \io_slave_araddr[24] ;
wire \io_slave_araddr[25] ;
wire \io_slave_araddr[26] ;
wire \io_slave_araddr[27] ;
wire \io_slave_araddr[28] ;
wire \io_slave_araddr[29] ;
wire \io_slave_araddr[30] ;
wire \io_slave_araddr[31] ;
wire \io_slave_arid[0] ;
wire \io_slave_arid[1] ;
wire \io_slave_arid[2] ;
wire \io_slave_arid[3] ;
wire \io_slave_arlen[0] ;
wire \io_slave_arlen[1] ;
wire \io_slave_arlen[2] ;
wire \io_slave_arlen[3] ;
wire \io_slave_arlen[4] ;
wire \io_slave_arlen[5] ;
wire \io_slave_arlen[6] ;
wire \io_slave_arlen[7] ;
wire \io_slave_arsize[0] ;
wire \io_slave_arsize[1] ;
wire \io_slave_arsize[2] ;
wire \io_slave_arburst[0] ;
wire \io_slave_arburst[1] ;
wire \io_slave_rresp[0] ;
wire \io_slave_rresp[1] ;
wire \io_slave_rdata[0] ;
wire \io_slave_rdata[1] ;
wire \io_slave_rdata[2] ;
wire \io_slave_rdata[3] ;
wire \io_slave_rdata[4] ;
wire \io_slave_rdata[5] ;
wire \io_slave_rdata[6] ;
wire \io_slave_rdata[7] ;
wire \io_slave_rdata[8] ;
wire \io_slave_rdata[9] ;
wire \io_slave_rdata[10] ;
wire \io_slave_rdata[11] ;
wire \io_slave_rdata[12] ;
wire \io_slave_rdata[13] ;
wire \io_slave_rdata[14] ;
wire \io_slave_rdata[15] ;
wire \io_slave_rdata[16] ;
wire \io_slave_rdata[17] ;
wire \io_slave_rdata[18] ;
wire \io_slave_rdata[19] ;
wire \io_slave_rdata[20] ;
wire \io_slave_rdata[21] ;
wire \io_slave_rdata[22] ;
wire \io_slave_rdata[23] ;
wire \io_slave_rdata[24] ;
wire \io_slave_rdata[25] ;
wire \io_slave_rdata[26] ;
wire \io_slave_rdata[27] ;
wire \io_slave_rdata[28] ;
wire \io_slave_rdata[29] ;
wire \io_slave_rdata[30] ;
wire \io_slave_rdata[31] ;
wire \io_slave_rid[0] ;
wire \io_slave_rid[1] ;
wire \io_slave_rid[2] ;
wire \io_slave_rid[3] ;
wire \ac_data[0] ;
wire \ac_data[1] ;
wire \ac_data[2] ;
wire \ac_data[3] ;
wire \ac_data[4] ;
wire \ac_data[5] ;
wire \ac_data[6] ;
wire \ac_data[7] ;
wire \ac_data[8] ;
wire \ac_data[9] ;
wire \ac_data[10] ;
wire \ac_data[11] ;
wire \ac_data[12] ;
wire \ac_data[13] ;
wire \ac_data[14] ;
wire \ac_data[15] ;
wire \ac_data[16] ;
wire \ac_data[17] ;
wire \ac_data[18] ;
wire \ac_data[19] ;
wire \ac_data[20] ;
wire \ac_data[21] ;
wire \ac_data[22] ;
wire \ac_data[23] ;
wire \ac_data[24] ;
wire \ac_data[25] ;
wire \ac_data[26] ;
wire \ac_data[27] ;
wire \ac_data[28] ;
wire \ac_data[29] ;
wire \ac_data[30] ;
wire \ac_data[31] ;
wire \al_wdata[0] ;
wire \al_wdata[1] ;
wire \al_wdata[2] ;
wire \al_wdata[3] ;
wire \al_wdata[4] ;
wire \al_wdata[5] ;
wire \al_wdata[6] ;
wire \al_wdata[7] ;
wire \al_wdata[8] ;
wire \al_wdata[9] ;
wire \al_wdata[10] ;
wire \al_wdata[11] ;
wire \al_wdata[12] ;
wire \al_wdata[13] ;
wire \al_wdata[14] ;
wire \al_wdata[15] ;
wire \al_wdata[16] ;
wire \al_wdata[17] ;
wire \al_wdata[18] ;
wire \al_wdata[19] ;
wire \al_wdata[20] ;
wire \al_wdata[21] ;
wire \al_wdata[22] ;
wire \al_wdata[23] ;
wire \al_wdata[24] ;
wire \al_wdata[25] ;
wire \al_wdata[26] ;
wire \al_wdata[27] ;
wire \al_wdata[28] ;
wire \al_wdata[29] ;
wire \al_wdata[30] ;
wire \al_wdata[31] ;
wire \al_wmask[0] ;
wire \al_wmask[1] ;
wire \ar_data[0] ;
wire \ar_data[1] ;
wire \ar_data[2] ;
wire \ar_data[3] ;
wire \ar_data[4] ;
wire \ar_data[5] ;
wire \ar_data[6] ;
wire \ar_data[7] ;
wire \ar_data[8] ;
wire \ar_data[9] ;
wire \ar_data[10] ;
wire \ar_data[11] ;
wire \ar_data[12] ;
wire \ar_data[13] ;
wire \ar_data[14] ;
wire \ar_data[15] ;
wire \ar_data[16] ;
wire \ar_data[17] ;
wire \ar_data[18] ;
wire \ar_data[19] ;
wire \ar_data[20] ;
wire \ar_data[21] ;
wire \ar_data[22] ;
wire \ar_data[23] ;
wire \ar_data[24] ;
wire \ar_data[25] ;
wire \ar_data[26] ;
wire \ar_data[27] ;
wire \ar_data[28] ;
wire \ar_data[29] ;
wire \ar_data[30] ;
wire \ar_data[31] ;
wire \ca_addr[0] ;
wire \ca_addr[1] ;
wire \ca_addr[2] ;
wire \ca_addr[3] ;
wire \ca_addr[4] ;
wire \ca_addr[5] ;
wire \ca_addr[6] ;
wire \ca_addr[7] ;
wire \ca_addr[8] ;
wire \ca_addr[9] ;
wire \ca_addr[10] ;
wire \ca_addr[11] ;
wire \ca_addr[12] ;
wire \ca_addr[13] ;
wire \ca_addr[14] ;
wire \ca_addr[15] ;
wire \ca_addr[16] ;
wire \ca_addr[17] ;
wire \ca_addr[18] ;
wire \ca_addr[19] ;
wire \ca_addr[20] ;
wire \ca_addr[21] ;
wire \ca_addr[22] ;
wire \ca_addr[23] ;
wire \ca_addr[24] ;
wire \ca_addr[25] ;
wire \ca_addr[26] ;
wire \ca_addr[27] ;
wire \ca_addr[28] ;
wire \ca_addr[29] ;
wire \ca_addr[30] ;
wire \ca_addr[31] ;
wire \cf_inst[0] ;
wire \cf_inst[1] ;
wire \cf_inst[2] ;
wire \cf_inst[3] ;
wire \cf_inst[4] ;
wire \cf_inst[5] ;
wire \cf_inst[6] ;
wire \cf_inst[7] ;
wire \cf_inst[8] ;
wire \cf_inst[9] ;
wire \cf_inst[10] ;
wire \cf_inst[11] ;
wire \cf_inst[12] ;
wire \cf_inst[13] ;
wire \cf_inst[14] ;
wire \cf_inst[15] ;
wire \cf_inst[16] ;
wire \cf_inst[17] ;
wire \cf_inst[18] ;
wire \cf_inst[19] ;
wire \cf_inst[20] ;
wire \cf_inst[21] ;
wire \cf_inst[22] ;
wire \cf_inst[23] ;
wire \cf_inst[24] ;
wire \cf_inst[25] ;
wire \cf_inst[26] ;
wire \cf_inst[27] ;
wire \cf_inst[28] ;
wire \cf_inst[29] ;
wire \cf_inst[30] ;
wire \cf_inst[31] ;
wire \de_pc[0] ;
wire \de_pc[1] ;
wire \de_pc[2] ;
wire \de_pc[3] ;
wire \de_pc[4] ;
wire \de_pc[5] ;
wire \de_pc[6] ;
wire \de_pc[7] ;
wire \de_pc[8] ;
wire \de_pc[9] ;
wire \de_pc[10] ;
wire \de_pc[11] ;
wire \de_pc[12] ;
wire \de_pc[13] ;
wire \de_pc[14] ;
wire \de_pc[15] ;
wire \de_pc[16] ;
wire \de_pc[17] ;
wire \de_pc[18] ;
wire \de_pc[19] ;
wire \de_pc[20] ;
wire \de_pc[21] ;
wire \de_pc[22] ;
wire \de_pc[23] ;
wire \de_pc[24] ;
wire \de_pc[25] ;
wire \de_pc[26] ;
wire \de_pc[27] ;
wire \de_pc[28] ;
wire \de_pc[29] ;
wire \de_pc[30] ;
wire \de_pc[31] ;
wire \ea_addr[0] ;
wire \ea_addr[1] ;
wire \ea_addr[2] ;
wire \ea_addr[3] ;
wire \ea_addr[4] ;
wire \ea_addr[5] ;
wire \ea_addr[6] ;
wire \ea_addr[7] ;
wire \ea_addr[8] ;
wire \ea_addr[9] ;
wire \ea_addr[10] ;
wire \ea_addr[11] ;
wire \ea_addr[12] ;
wire \ea_addr[13] ;
wire \ea_addr[14] ;
wire \ea_addr[15] ;
wire \ea_addr[16] ;
wire \ea_addr[17] ;
wire \ea_addr[18] ;
wire \ea_addr[19] ;
wire \ea_addr[20] ;
wire \ea_addr[21] ;
wire \ea_addr[22] ;
wire \ea_addr[23] ;
wire \ea_addr[24] ;
wire \ea_addr[25] ;
wire \ea_addr[26] ;
wire \ea_addr[27] ;
wire \ea_addr[28] ;
wire \ea_addr[29] ;
wire \ea_addr[30] ;
wire \ea_addr[31] ;
wire \ea_ard[0] ;
wire \ea_ard[1] ;
wire \ea_ard[2] ;
wire \ea_ard[3] ;
wire \ea_errtp[0] ;
wire \ea_mask[0] ;
wire \ea_mask[1] ;
wire \ea_pc[0] ;
wire \ea_pc[1] ;
wire \ea_pc[2] ;
wire \ea_pc[3] ;
wire \ea_pc[4] ;
wire \ea_pc[5] ;
wire \ea_pc[6] ;
wire \ea_pc[7] ;
wire \ea_pc[8] ;
wire \ea_pc[9] ;
wire \ea_pc[10] ;
wire \ea_pc[11] ;
wire \ea_pc[12] ;
wire \ea_pc[13] ;
wire \ea_pc[14] ;
wire \ea_pc[15] ;
wire \ea_pc[16] ;
wire \ea_pc[17] ;
wire \ea_pc[18] ;
wire \ea_pc[19] ;
wire \ea_pc[20] ;
wire \ea_pc[21] ;
wire \ea_pc[22] ;
wire \ea_pc[23] ;
wire \ea_pc[24] ;
wire \ea_pc[25] ;
wire \ea_pc[26] ;
wire \ea_pc[27] ;
wire \ea_pc[28] ;
wire \ea_pc[29] ;
wire \ea_pc[30] ;
wire \ea_pc[31] ;
wire \ea_wdata[0] ;
wire \ea_wdata[1] ;
wire \ea_wdata[2] ;
wire \ea_wdata[3] ;
wire \ea_wdata[4] ;
wire \ea_wdata[5] ;
wire \ea_wdata[6] ;
wire \ea_wdata[7] ;
wire \ea_wdata[8] ;
wire \ea_wdata[9] ;
wire \ea_wdata[10] ;
wire \ea_wdata[11] ;
wire \ea_wdata[12] ;
wire \ea_wdata[13] ;
wire \ea_wdata[14] ;
wire \ea_wdata[15] ;
wire \ea_wdata[16] ;
wire \ea_wdata[17] ;
wire \ea_wdata[18] ;
wire \ea_wdata[19] ;
wire \ea_wdata[20] ;
wire \ea_wdata[21] ;
wire \ea_wdata[22] ;
wire \ea_wdata[23] ;
wire \ea_wdata[24] ;
wire \ea_wdata[25] ;
wire \ea_wdata[26] ;
wire \ea_wdata[27] ;
wire \ea_wdata[28] ;
wire \ea_wdata[29] ;
wire \ea_wdata[30] ;
wire \ea_wdata[31] ;
wire \fc_addr[0] ;
wire \fc_addr[1] ;
wire \fc_addr[2] ;
wire \fc_addr[3] ;
wire \fc_addr[4] ;
wire \fc_addr[5] ;
wire \fc_addr[6] ;
wire \fc_addr[7] ;
wire \fc_addr[8] ;
wire \fc_addr[9] ;
wire \fc_addr[10] ;
wire \fc_addr[11] ;
wire \fc_addr[12] ;
wire \fc_addr[13] ;
wire \fc_addr[14] ;
wire \fc_addr[15] ;
wire \fc_addr[16] ;
wire \fc_addr[17] ;
wire \fc_addr[18] ;
wire \fc_addr[19] ;
wire \fc_addr[20] ;
wire \fc_addr[21] ;
wire \fc_addr[22] ;
wire \fc_addr[23] ;
wire \fc_addr[24] ;
wire \fc_addr[25] ;
wire \fc_addr[26] ;
wire \fc_addr[27] ;
wire \fc_addr[28] ;
wire \fc_addr[29] ;
wire \fc_addr[30] ;
wire \fc_addr[31] ;
wire \fd_inst[0] ;
wire \fd_inst[1] ;
wire \fd_inst[2] ;
wire \fd_inst[3] ;
wire \fd_inst[4] ;
wire \fd_inst[5] ;
wire \fd_inst[6] ;
wire \fd_inst[7] ;
wire \fd_inst[8] ;
wire \fd_inst[9] ;
wire \fd_inst[10] ;
wire \fd_inst[11] ;
wire \fd_inst[12] ;
wire \fd_inst[13] ;
wire \fd_inst[14] ;
wire \fd_inst[15] ;
wire \fd_inst[16] ;
wire \fd_inst[17] ;
wire \fd_inst[18] ;
wire \fd_inst[19] ;
wire \fd_inst[20] ;
wire \fd_inst[21] ;
wire \fd_inst[22] ;
wire \fd_inst[23] ;
wire \fd_inst[24] ;
wire \fd_inst[25] ;
wire \fd_inst[26] ;
wire \fd_inst[27] ;
wire \fd_inst[28] ;
wire \fd_inst[29] ;
wire \fd_inst[30] ;
wire \fd_inst[31] ;
wire \u_arbiter.raddr[0] ;
wire \u_arbiter.raddr[1] ;
wire \u_arbiter.raddr[2] ;
wire \u_arbiter.raddr[3] ;
wire \u_arbiter.raddr[4] ;
wire \u_arbiter.raddr[5] ;
wire \u_arbiter.raddr[6] ;
wire \u_arbiter.raddr[7] ;
wire \u_arbiter.raddr[8] ;
wire \u_arbiter.raddr[9] ;
wire \u_arbiter.raddr[10] ;
wire \u_arbiter.raddr[11] ;
wire \u_arbiter.raddr[12] ;
wire \u_arbiter.raddr[13] ;
wire \u_arbiter.raddr[14] ;
wire \u_arbiter.raddr[15] ;
wire \u_arbiter.raddr[16] ;
wire \u_arbiter.raddr[17] ;
wire \u_arbiter.raddr[18] ;
wire \u_arbiter.raddr[19] ;
wire \u_arbiter.raddr[20] ;
wire \u_arbiter.raddr[21] ;
wire \u_arbiter.raddr[22] ;
wire \u_arbiter.raddr[23] ;
wire \u_arbiter.raddr[24] ;
wire \u_arbiter.raddr[25] ;
wire \u_arbiter.raddr[26] ;
wire \u_arbiter.raddr[27] ;
wire \u_arbiter.raddr[28] ;
wire \u_arbiter.raddr[29] ;
wire \u_arbiter.raddr[30] ;
wire \u_arbiter.raddr[31] ;
wire \u_arbiter.rmask[0] ;
wire \u_arbiter.rmask[1] ;
wire \u_arbiter.wbaddr[0] ;
wire \u_arbiter.wbaddr[1] ;
wire \u_arbiter.wbaddr[2] ;
wire \u_arbiter.wbaddr[3] ;
wire \u_exu.acsrd[0] ;
wire \u_exu.acsrd[1] ;
wire \u_exu.acsrd[2] ;
wire \u_exu.acsrd[3] ;
wire \u_exu.acsrd[4] ;
wire \u_exu.acsrd[5] ;
wire \u_exu.acsrd[6] ;
wire \u_exu.acsrd[7] ;
wire \u_exu.acsrd[8] ;
wire \u_exu.acsrd[9] ;
wire \u_exu.acsrd[10] ;
wire \u_exu.acsrd[11] ;
wire \u_exu.alu_ctrl[0] ;
wire \u_exu.alu_ctrl[1] ;
wire \u_exu.alu_ctrl[2] ;
wire \u_exu.alu_ctrl[3] ;
wire \u_exu.alu_ctrl[4] ;
wire \u_exu.alu_ctrl[5] ;
wire \u_exu.alu_ctrl[6] ;
wire \u_exu.alu_p1[0] ;
wire \u_exu.alu_p1[1] ;
wire \u_exu.alu_p1[2] ;
wire \u_exu.alu_p1[3] ;
wire \u_exu.alu_p1[4] ;
wire \u_exu.alu_p1[5] ;
wire \u_exu.alu_p1[6] ;
wire \u_exu.alu_p1[7] ;
wire \u_exu.alu_p1[8] ;
wire \u_exu.alu_p1[9] ;
wire \u_exu.alu_p1[10] ;
wire \u_exu.alu_p1[11] ;
wire \u_exu.alu_p1[12] ;
wire \u_exu.alu_p1[13] ;
wire \u_exu.alu_p1[14] ;
wire \u_exu.alu_p1[15] ;
wire \u_exu.alu_p1[16] ;
wire \u_exu.alu_p1[17] ;
wire \u_exu.alu_p1[18] ;
wire \u_exu.alu_p1[19] ;
wire \u_exu.alu_p1[20] ;
wire \u_exu.alu_p1[21] ;
wire \u_exu.alu_p1[22] ;
wire \u_exu.alu_p1[23] ;
wire \u_exu.alu_p1[24] ;
wire \u_exu.alu_p1[25] ;
wire \u_exu.alu_p1[26] ;
wire \u_exu.alu_p1[27] ;
wire \u_exu.alu_p1[28] ;
wire \u_exu.alu_p1[29] ;
wire \u_exu.alu_p1[30] ;
wire \u_exu.alu_p1[31] ;
wire \u_exu.alu_p2[0] ;
wire \u_exu.alu_p2[1] ;
wire \u_exu.alu_p2[2] ;
wire \u_exu.alu_p2[3] ;
wire \u_exu.alu_p2[4] ;
wire \u_exu.alu_p2[5] ;
wire \u_exu.alu_p2[6] ;
wire \u_exu.alu_p2[7] ;
wire \u_exu.alu_p2[8] ;
wire \u_exu.alu_p2[9] ;
wire \u_exu.alu_p2[10] ;
wire \u_exu.alu_p2[11] ;
wire \u_exu.alu_p2[12] ;
wire \u_exu.alu_p2[13] ;
wire \u_exu.alu_p2[14] ;
wire \u_exu.alu_p2[15] ;
wire \u_exu.alu_p2[16] ;
wire \u_exu.alu_p2[17] ;
wire \u_exu.alu_p2[18] ;
wire \u_exu.alu_p2[19] ;
wire \u_exu.alu_p2[20] ;
wire \u_exu.alu_p2[21] ;
wire \u_exu.alu_p2[22] ;
wire \u_exu.alu_p2[23] ;
wire \u_exu.alu_p2[24] ;
wire \u_exu.alu_p2[25] ;
wire \u_exu.alu_p2[26] ;
wire \u_exu.alu_p2[27] ;
wire \u_exu.alu_p2[28] ;
wire \u_exu.alu_p2[29] ;
wire \u_exu.alu_p2[30] ;
wire \u_exu.alu_p2[31] ;
wire \u_exu.ecsr[0] ;
wire \u_exu.ecsr[1] ;
wire \u_exu.ecsr[2] ;
wire \u_exu.ecsr[3] ;
wire \u_exu.ecsr[4] ;
wire \u_exu.ecsr[5] ;
wire \u_exu.ecsr[6] ;
wire \u_exu.ecsr[7] ;
wire \u_exu.ecsr[8] ;
wire \u_exu.ecsr[9] ;
wire \u_exu.ecsr[10] ;
wire \u_exu.ecsr[11] ;
wire \u_exu.ecsr[12] ;
wire \u_exu.ecsr[13] ;
wire \u_exu.ecsr[14] ;
wire \u_exu.ecsr[15] ;
wire \u_exu.ecsr[16] ;
wire \u_exu.ecsr[17] ;
wire \u_exu.ecsr[18] ;
wire \u_exu.ecsr[19] ;
wire \u_exu.ecsr[20] ;
wire \u_exu.ecsr[21] ;
wire \u_exu.ecsr[22] ;
wire \u_exu.ecsr[23] ;
wire \u_exu.ecsr[24] ;
wire \u_exu.ecsr[25] ;
wire \u_exu.ecsr[26] ;
wire \u_exu.ecsr[27] ;
wire \u_exu.ecsr[28] ;
wire \u_exu.ecsr[29] ;
wire \u_exu.ecsr[30] ;
wire \u_exu.ecsr[31] ;
wire \u_exu.eopt[0] ;
wire \u_exu.eopt[1] ;
wire \u_exu.eopt[2] ;
wire \u_exu.eopt[3] ;
wire \u_exu.eopt[4] ;
wire \u_exu.eopt[5] ;
wire \u_exu.eopt[6] ;
wire \u_exu.eopt[7] ;
wire \u_exu.eopt[8] ;
wire \u_exu.eopt[9] ;
wire \u_exu.eopt[10] ;
wire \u_exu.eopt[11] ;
wire \u_exu.eopt[12] ;
wire \u_exu.eopt[13] ;
wire \u_exu.eopt[14] ;
wire \u_exu.eopt[15] ;
wire \u_exu.rlock[0] ;
wire \u_exu.rlock[1] ;
wire \u_exu.rlock[2] ;
wire \u_exu.rlock[3] ;
wire \u_exu.rlock[4] ;
wire \u_exu.rlock[5] ;
wire \u_exu.rlock[6] ;
wire \u_exu.rlock[7] ;
wire \u_exu.rlock[8] ;
wire \u_exu.rlock[9] ;
wire \u_exu.rlock[10] ;
wire \u_exu.rlock[11] ;
wire \u_exu.rlock[12] ;
wire \u_exu.rlock[13] ;
wire \u_exu.rlock[14] ;
wire \u_exu.rlock[15] ;
wire \u_icache.count[0] ;
wire \u_icache.count[1] ;
wire \u_icache.count[2] ;
wire \u_icache.cvalids[0] ;
wire \u_icache.cvalids[1] ;
wire \u_idu.imm_auipc_lui[0] ;
wire \u_idu.imm_auipc_lui[1] ;
wire \u_idu.imm_auipc_lui[2] ;
wire \u_idu.imm_auipc_lui[3] ;
wire \u_idu.imm_auipc_lui[4] ;
wire \u_idu.imm_auipc_lui[5] ;
wire \u_idu.imm_auipc_lui[6] ;
wire \u_idu.imm_auipc_lui[7] ;
wire \u_idu.imm_auipc_lui[8] ;
wire \u_idu.imm_auipc_lui[9] ;
wire \u_idu.imm_auipc_lui[10] ;
wire \u_idu.imm_auipc_lui[11] ;
wire \u_idu.imm_auipc_lui[12] ;
wire \u_idu.imm_auipc_lui[13] ;
wire \u_idu.imm_auipc_lui[14] ;
wire \u_idu.imm_auipc_lui[15] ;
wire \u_idu.imm_auipc_lui[16] ;
wire \u_idu.imm_auipc_lui[17] ;
wire \u_idu.imm_auipc_lui[18] ;
wire \u_idu.imm_auipc_lui[19] ;
wire \u_idu.imm_auipc_lui[20] ;
wire \u_idu.imm_auipc_lui[21] ;
wire \u_idu.imm_auipc_lui[22] ;
wire \u_idu.imm_auipc_lui[23] ;
wire \u_idu.imm_auipc_lui[24] ;
wire \u_idu.imm_auipc_lui[25] ;
wire \u_idu.imm_auipc_lui[26] ;
wire \u_idu.imm_auipc_lui[27] ;
wire \u_idu.imm_auipc_lui[28] ;
wire \u_idu.imm_auipc_lui[29] ;
wire \u_idu.imm_auipc_lui[30] ;
wire \u_idu.imm_auipc_lui[31] ;
wire \u_idu.imm_branch[0] ;
wire \u_idu.imm_branch[1] ;
wire \u_idu.imm_branch[2] ;
wire \u_idu.imm_branch[3] ;
wire \u_idu.imm_branch[4] ;
wire \u_idu.imm_branch[5] ;
wire \u_idu.imm_branch[6] ;
wire \u_idu.imm_branch[7] ;
wire \u_idu.imm_branch[8] ;
wire \u_idu.imm_branch[9] ;
wire \u_idu.imm_branch[10] ;
wire \u_idu.imm_branch[11] ;
wire \u_idu.inst[0] ;
wire \u_idu.inst[1] ;
wire \u_idu.inst[2] ;
wire \u_idu.inst[3] ;
wire \u_idu.inst[4] ;
wire \u_idu.inst[5] ;
wire \u_idu.inst[6] ;
wire \u_lsu.rcount[0] ;
wire \u_lsu.rcount[1] ;
wire \u_lsu.rcount[2] ;
wire \u_lsu.rcount[3] ;
wire \u_lsu.rcount[4] ;
wire \u_lsu.rcount[5] ;
wire \u_lsu.rcount[6] ;
wire \u_lsu.rcount[7] ;
wire \u_lsu.u_clint.mtime[0] ;
wire \u_lsu.u_clint.mtime[1] ;
wire \u_lsu.u_clint.mtime[2] ;
wire \u_lsu.u_clint.mtime[3] ;
wire \u_lsu.u_clint.mtime[4] ;
wire \u_lsu.u_clint.mtime[5] ;
wire \u_lsu.u_clint.mtime[6] ;
wire \u_lsu.u_clint.mtime[7] ;
wire \u_lsu.u_clint.mtime[8] ;
wire \u_lsu.u_clint.mtime[9] ;
wire \u_lsu.u_clint.mtime[10] ;
wire \u_lsu.u_clint.mtime[11] ;
wire \u_lsu.u_clint.mtime[12] ;
wire \u_lsu.u_clint.mtime[13] ;
wire \u_lsu.u_clint.mtime[14] ;
wire \u_lsu.u_clint.mtime[15] ;
wire \u_lsu.u_clint.mtime[16] ;
wire \u_lsu.u_clint.mtime[17] ;
wire \u_lsu.u_clint.mtime[18] ;
wire \u_lsu.u_clint.mtime[19] ;
wire \u_lsu.u_clint.mtime[20] ;
wire \u_lsu.u_clint.mtime[21] ;
wire \u_lsu.u_clint.mtime[22] ;
wire \u_lsu.u_clint.mtime[23] ;
wire \u_lsu.u_clint.mtime[24] ;
wire \u_lsu.u_clint.mtime[25] ;
wire \u_lsu.u_clint.mtime[26] ;
wire \u_lsu.u_clint.mtime[27] ;
wire \u_lsu.u_clint.mtime[28] ;
wire \u_lsu.u_clint.mtime[29] ;
wire \u_lsu.u_clint.mtime[30] ;
wire \u_lsu.u_clint.mtime[31] ;
wire \u_lsu.u_clint.mtime[32] ;
wire \u_lsu.u_clint.mtime[33] ;
wire \u_lsu.u_clint.mtime[34] ;
wire \u_lsu.u_clint.mtime[35] ;
wire \u_lsu.u_clint.mtime[36] ;
wire \u_lsu.u_clint.mtime[37] ;
wire \u_lsu.u_clint.mtime[38] ;
wire \u_lsu.u_clint.mtime[39] ;
wire \u_lsu.u_clint.mtime[40] ;
wire \u_lsu.u_clint.mtime[41] ;
wire \u_lsu.u_clint.mtime[42] ;
wire \u_lsu.u_clint.mtime[43] ;
wire \u_lsu.u_clint.mtime[44] ;
wire \u_lsu.u_clint.mtime[45] ;
wire \u_lsu.u_clint.mtime[46] ;
wire \u_lsu.u_clint.mtime[47] ;
wire \u_lsu.u_clint.mtime[48] ;
wire \u_lsu.u_clint.mtime[49] ;
wire \u_lsu.u_clint.mtime[50] ;
wire \u_lsu.u_clint.mtime[51] ;
wire \u_lsu.u_clint.mtime[52] ;
wire \u_lsu.u_clint.mtime[53] ;
wire \u_lsu.u_clint.mtime[54] ;
wire \u_lsu.u_clint.mtime[55] ;
wire \u_lsu.u_clint.mtime[56] ;
wire \u_lsu.u_clint.mtime[57] ;
wire \u_lsu.u_clint.mtime[58] ;
wire \u_lsu.u_clint.mtime[59] ;
wire \u_lsu.u_clint.mtime[60] ;
wire \u_lsu.u_clint.mtime[61] ;
wire \u_lsu.u_clint.mtime[62] ;
wire \u_lsu.u_clint.mtime[63] ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D[0] ;

assign io_master_wlast = io_master_wvalid ;
assign io_master_awaddr[0] = \io_master_awaddr[0] ;
assign io_master_awaddr[1] = \io_master_awaddr[1] ;
assign io_master_awaddr[2] = \io_master_awaddr[2] ;
assign io_master_awaddr[3] = \io_master_awaddr[3] ;
assign io_master_awaddr[4] = \io_master_awaddr[4] ;
assign io_master_awaddr[5] = \io_master_awaddr[5] ;
assign io_master_awaddr[6] = \io_master_awaddr[6] ;
assign io_master_awaddr[7] = \io_master_awaddr[7] ;
assign io_master_awaddr[8] = \io_master_awaddr[8] ;
assign io_master_awaddr[9] = \io_master_awaddr[9] ;
assign io_master_awaddr[10] = \io_master_awaddr[10] ;
assign io_master_awaddr[11] = \io_master_awaddr[11] ;
assign io_master_awaddr[12] = \io_master_awaddr[12] ;
assign io_master_awaddr[13] = \io_master_awaddr[13] ;
assign io_master_awaddr[14] = \io_master_awaddr[14] ;
assign io_master_awaddr[15] = \io_master_awaddr[15] ;
assign io_master_awaddr[16] = \io_master_awaddr[16] ;
assign io_master_awaddr[17] = \io_master_awaddr[17] ;
assign io_master_awaddr[18] = \io_master_awaddr[18] ;
assign io_master_awaddr[19] = \io_master_awaddr[19] ;
assign io_master_awaddr[20] = \io_master_awaddr[20] ;
assign io_master_awaddr[21] = \io_master_awaddr[21] ;
assign io_master_awaddr[22] = \io_master_awaddr[22] ;
assign io_master_awaddr[23] = \io_master_awaddr[23] ;
assign io_master_awaddr[24] = \io_master_awaddr[24] ;
assign io_master_awaddr[25] = \io_master_awaddr[25] ;
assign io_master_awaddr[26] = \io_master_awaddr[26] ;
assign io_master_awaddr[27] = \io_master_awaddr[27] ;
assign io_master_awaddr[28] = \io_master_awaddr[28] ;
assign io_master_awaddr[29] = \io_master_awaddr[29] ;
assign io_master_awaddr[30] = \io_master_awaddr[30] ;
assign io_master_awaddr[31] = \io_master_awaddr[31] ;
assign io_master_arburst[1] = \io_master_awid[0] ;
assign io_master_arburst[1] = \io_master_awid[1] ;
assign io_master_arburst[1] = \io_master_awid[2] ;
assign io_master_arburst[1] = \io_master_awid[3] ;
assign io_master_arburst[1] = \io_master_awlen[0] ;
assign io_master_arburst[1] = \io_master_awlen[1] ;
assign io_master_arburst[1] = \io_master_awlen[2] ;
assign io_master_arburst[1] = \io_master_awlen[3] ;
assign io_master_arburst[1] = \io_master_awlen[4] ;
assign io_master_arburst[1] = \io_master_awlen[5] ;
assign io_master_arburst[1] = \io_master_awlen[6] ;
assign io_master_arburst[1] = \io_master_awlen[7] ;
assign io_master_awsize[0] = \io_master_awsize[0] ;
assign io_master_awsize[1] = \io_master_awsize[1] ;
assign io_master_arburst[1] = \io_master_awsize[2] ;
assign io_master_arburst[1] = \io_master_awburst[0] ;
assign io_master_arburst[1] = \io_master_awburst[1] ;
assign io_master_wdata[0] = \io_master_wdata[0] ;
assign io_master_wdata[1] = \io_master_wdata[1] ;
assign io_master_wdata[2] = \io_master_wdata[2] ;
assign io_master_wdata[3] = \io_master_wdata[3] ;
assign io_master_wdata[4] = \io_master_wdata[4] ;
assign io_master_wdata[5] = \io_master_wdata[5] ;
assign io_master_wdata[6] = \io_master_wdata[6] ;
assign io_master_wdata[7] = \io_master_wdata[7] ;
assign io_master_wdata[8] = \io_master_wdata[8] ;
assign io_master_wdata[9] = \io_master_wdata[9] ;
assign io_master_wdata[10] = \io_master_wdata[10] ;
assign io_master_wdata[11] = \io_master_wdata[11] ;
assign io_master_wdata[12] = \io_master_wdata[12] ;
assign io_master_wdata[13] = \io_master_wdata[13] ;
assign io_master_wdata[14] = \io_master_wdata[14] ;
assign io_master_wdata[15] = \io_master_wdata[15] ;
assign io_master_wdata[16] = \io_master_wdata[16] ;
assign io_master_wdata[17] = \io_master_wdata[17] ;
assign io_master_wdata[18] = \io_master_wdata[18] ;
assign io_master_wdata[19] = \io_master_wdata[19] ;
assign io_master_wdata[20] = \io_master_wdata[20] ;
assign io_master_wdata[21] = \io_master_wdata[21] ;
assign io_master_wdata[22] = \io_master_wdata[22] ;
assign io_master_wdata[23] = \io_master_wdata[23] ;
assign io_master_wdata[24] = \io_master_wdata[24] ;
assign io_master_wdata[25] = \io_master_wdata[25] ;
assign io_master_wdata[26] = \io_master_wdata[26] ;
assign io_master_wdata[27] = \io_master_wdata[27] ;
assign io_master_wdata[28] = \io_master_wdata[28] ;
assign io_master_wdata[29] = \io_master_wdata[29] ;
assign io_master_wdata[30] = \io_master_wdata[30] ;
assign io_master_wdata[31] = \io_master_wdata[31] ;
assign io_master_wstrb[0] = \io_master_wstrb[0] ;
assign io_master_wstrb[1] = \io_master_wstrb[1] ;
assign io_master_wstrb[2] = \io_master_wstrb[2] ;
assign io_master_wstrb[3] = \io_master_wstrb[3] ;
assign io_master_araddr[0] = \io_master_araddr[0] ;
assign io_master_araddr[1] = \io_master_araddr[1] ;
assign io_master_araddr[2] = \io_master_araddr[2] ;
assign io_master_araddr[3] = \io_master_araddr[3] ;
assign io_master_araddr[4] = \io_master_araddr[4] ;
assign io_master_araddr[5] = \io_master_araddr[5] ;
assign io_master_araddr[6] = \io_master_araddr[6] ;
assign io_master_araddr[7] = \io_master_araddr[7] ;
assign io_master_araddr[8] = \io_master_araddr[8] ;
assign io_master_araddr[9] = \io_master_araddr[9] ;
assign io_master_araddr[10] = \io_master_araddr[10] ;
assign io_master_araddr[11] = \io_master_araddr[11] ;
assign io_master_araddr[12] = \io_master_araddr[12] ;
assign io_master_araddr[13] = \io_master_araddr[13] ;
assign io_master_araddr[14] = \io_master_araddr[14] ;
assign io_master_araddr[15] = \io_master_araddr[15] ;
assign io_master_araddr[16] = \io_master_araddr[16] ;
assign io_master_araddr[17] = \io_master_araddr[17] ;
assign io_master_araddr[18] = \io_master_araddr[18] ;
assign io_master_araddr[19] = \io_master_araddr[19] ;
assign io_master_araddr[20] = \io_master_araddr[20] ;
assign io_master_araddr[21] = \io_master_araddr[21] ;
assign io_master_araddr[22] = \io_master_araddr[22] ;
assign io_master_araddr[23] = \io_master_araddr[23] ;
assign io_master_araddr[24] = \io_master_araddr[24] ;
assign io_master_araddr[25] = \io_master_araddr[25] ;
assign io_master_araddr[26] = \io_master_araddr[26] ;
assign io_master_araddr[27] = \io_master_araddr[27] ;
assign io_master_araddr[28] = \io_master_araddr[28] ;
assign io_master_araddr[29] = \io_master_araddr[29] ;
assign io_master_araddr[30] = \io_master_araddr[30] ;
assign io_master_araddr[31] = \io_master_araddr[31] ;
assign io_master_arburst[1] = \io_master_arid[0] ;
assign io_master_arburst[1] = \io_master_arid[1] ;
assign io_master_arburst[1] = \io_master_arid[2] ;
assign io_master_arburst[1] = \io_master_arid[3] ;
assign io_master_arburst[0] = \io_master_arlen[0] ;
assign io_master_arburst[0] = \io_master_arlen[1] ;
assign io_master_arburst[1] = \io_master_arlen[2] ;
assign io_master_arburst[1] = \io_master_arlen[3] ;
assign io_master_arburst[1] = \io_master_arlen[4] ;
assign io_master_arburst[1] = \io_master_arlen[5] ;
assign io_master_arburst[1] = \io_master_arlen[6] ;
assign io_master_arburst[1] = \io_master_arlen[7] ;
assign io_master_arsize[0] = \io_master_arsize[0] ;
assign io_master_arsize[1] = \io_master_arsize[1] ;
assign io_master_arburst[1] = \io_master_arsize[2] ;
assign io_master_arburst[0] = \io_master_arburst[0] ;
assign io_master_arburst[1] = \io_master_arburst[1] ;
assign \io_master_rdata[0] = io_master_rdata[0] ;
assign \io_master_rdata[1] = io_master_rdata[1] ;
assign \io_master_rdata[2] = io_master_rdata[2] ;
assign \io_master_rdata[3] = io_master_rdata[3] ;
assign \io_master_rdata[4] = io_master_rdata[4] ;
assign \io_master_rdata[5] = io_master_rdata[5] ;
assign \io_master_rdata[6] = io_master_rdata[6] ;
assign \io_master_rdata[7] = io_master_rdata[7] ;
assign \io_master_rdata[8] = io_master_rdata[8] ;
assign \io_master_rdata[9] = io_master_rdata[9] ;
assign \io_master_rdata[10] = io_master_rdata[10] ;
assign \io_master_rdata[11] = io_master_rdata[11] ;
assign \io_master_rdata[12] = io_master_rdata[12] ;
assign \io_master_rdata[13] = io_master_rdata[13] ;
assign \io_master_rdata[14] = io_master_rdata[14] ;
assign \io_master_rdata[15] = io_master_rdata[15] ;
assign \io_master_rdata[16] = io_master_rdata[16] ;
assign \io_master_rdata[17] = io_master_rdata[17] ;
assign \io_master_rdata[18] = io_master_rdata[18] ;
assign \io_master_rdata[19] = io_master_rdata[19] ;
assign \io_master_rdata[20] = io_master_rdata[20] ;
assign \io_master_rdata[21] = io_master_rdata[21] ;
assign \io_master_rdata[22] = io_master_rdata[22] ;
assign \io_master_rdata[23] = io_master_rdata[23] ;
assign \io_master_rdata[24] = io_master_rdata[24] ;
assign \io_master_rdata[25] = io_master_rdata[25] ;
assign \io_master_rdata[26] = io_master_rdata[26] ;
assign \io_master_rdata[27] = io_master_rdata[27] ;
assign \io_master_rdata[28] = io_master_rdata[28] ;
assign \io_master_rdata[29] = io_master_rdata[29] ;
assign \io_master_rdata[30] = io_master_rdata[30] ;
assign \io_master_rdata[31] = io_master_rdata[31] ;

INV_X1 _07572_ ( .A(\ea_mask[1] ), .ZN(_00627_ ) );
INV_X1 _07573_ ( .A(\ea_mask[0] ), .ZN(_00628_ ) );
AOI21_X1 _07574_ ( .A(\u_exu.eopt[15] ), .B1(_00627_ ), .B2(_00628_ ), .ZN(_00629_ ) );
OR2_X1 _07575_ ( .A1(_00629_ ), .A2(fanout_net_5 ), .ZN(_00630_ ) );
AOI21_X1 _07576_ ( .A(\u_arbiter.working ), .B1(_00630_ ), .B2(icah_valid ), .ZN(_00631_ ) );
AND2_X2 _07577_ ( .A1(_00631_ ), .A2(exu_valid ), .ZN(_00632_ ) );
AND2_X1 _07578_ ( .A1(_00632_ ), .A2(fanout_net_5 ), .ZN(_00633_ ) );
BUF_X4 _07579_ ( .A(_00633_ ), .Z(_00634_ ) );
INV_X1 _07580_ ( .A(_00634_ ), .ZN(_00635_ ) );
BUF_X4 _07581_ ( .A(_00635_ ), .Z(_00636_ ) );
BUF_X4 _07582_ ( .A(_00636_ ), .Z(_00637_ ) );
NOR2_X1 _07583_ ( .A1(\u_idu.imm_auipc_lui[28] ), .A2(\u_idu.imm_auipc_lui[29] ), .ZN(_00638_ ) );
NOR2_X1 _07584_ ( .A1(\u_idu.imm_auipc_lui[27] ), .A2(\u_idu.imm_auipc_lui[26] ), .ZN(_00639_ ) );
AND2_X1 _07585_ ( .A1(_00638_ ), .A2(_00639_ ), .ZN(_00640_ ) );
NOR2_X1 _07586_ ( .A1(\u_idu.imm_auipc_lui[31] ), .A2(\u_idu.imm_auipc_lui[30] ), .ZN(_00641_ ) );
AND2_X1 _07587_ ( .A1(_00640_ ), .A2(_00641_ ), .ZN(_00642_ ) );
NOR2_X1 _07588_ ( .A1(\u_idu.imm_auipc_lui[14] ), .A2(\u_idu.imm_auipc_lui[25] ), .ZN(_00643_ ) );
AND3_X1 _07589_ ( .A1(_00642_ ), .A2(\u_idu.imm_auipc_lui[13] ), .A3(_00643_ ), .ZN(_00644_ ) );
INV_X1 _07590_ ( .A(\u_idu.imm_auipc_lui[12] ), .ZN(_00645_ ) );
AND3_X1 _07591_ ( .A1(_00641_ ), .A2(_00645_ ), .A3(\u_idu.imm_auipc_lui[13] ), .ZN(_00646_ ) );
INV_X1 _07592_ ( .A(\u_idu.imm_auipc_lui[14] ), .ZN(_00647_ ) );
NOR2_X1 _07593_ ( .A1(_00647_ ), .A2(\u_idu.imm_auipc_lui[25] ), .ZN(_00648_ ) );
AND3_X1 _07594_ ( .A1(_00646_ ), .A2(_00640_ ), .A3(_00648_ ), .ZN(_00649_ ) );
NOR2_X1 _07595_ ( .A1(_00644_ ), .A2(_00649_ ), .ZN(_00650_ ) );
NOR2_X1 _07596_ ( .A1(_00645_ ), .A2(\u_idu.imm_auipc_lui[13] ), .ZN(_00651_ ) );
AND3_X1 _07597_ ( .A1(_00640_ ), .A2(_00651_ ), .A3(_00648_ ), .ZN(_00652_ ) );
INV_X1 _07598_ ( .A(\u_idu.imm_auipc_lui[31] ), .ZN(_00653_ ) );
NAND2_X1 _07599_ ( .A1(_00652_ ), .A2(_00653_ ), .ZN(_00654_ ) );
NAND4_X1 _07600_ ( .A1(_00640_ ), .A2(_00651_ ), .A3(_00641_ ), .A4(_00643_ ), .ZN(_00655_ ) );
AND2_X1 _07601_ ( .A1(_00654_ ), .A2(_00655_ ), .ZN(_00656_ ) );
NOR2_X1 _07602_ ( .A1(\u_idu.imm_auipc_lui[12] ), .A2(\u_idu.imm_auipc_lui[13] ), .ZN(_00657_ ) );
AND3_X1 _07603_ ( .A1(_00640_ ), .A2(_00643_ ), .A3(_00657_ ), .ZN(_00658_ ) );
NAND2_X1 _07604_ ( .A1(_00658_ ), .A2(_00653_ ), .ZN(_00659_ ) );
AND2_X1 _07605_ ( .A1(\u_idu.imm_auipc_lui[12] ), .A2(\u_idu.imm_auipc_lui[13] ), .ZN(_00660_ ) );
OAI211_X1 _07606_ ( .A(_00642_ ), .B(_00648_ ), .C1(_00657_ ), .C2(_00660_ ), .ZN(_00661_ ) );
NAND4_X1 _07607_ ( .A1(_00650_ ), .A2(_00656_ ), .A3(_00659_ ), .A4(_00661_ ), .ZN(_00662_ ) );
AND2_X1 _07608_ ( .A1(\u_idu.inst[0] ), .A2(\u_idu.inst[1] ), .ZN(_00663_ ) );
NOR2_X1 _07609_ ( .A1(\u_idu.inst[3] ), .A2(\u_idu.inst[2] ), .ZN(_00664_ ) );
AND2_X2 _07610_ ( .A1(_00663_ ), .A2(_00664_ ), .ZN(_00665_ ) );
NAND2_X1 _07611_ ( .A1(\u_idu.inst[5] ), .A2(\u_idu.inst[4] ), .ZN(_00666_ ) );
NOR2_X1 _07612_ ( .A1(_00666_ ), .A2(\u_idu.inst[6] ), .ZN(_00667_ ) );
AND2_X2 _07613_ ( .A1(_00665_ ), .A2(_00667_ ), .ZN(_00668_ ) );
NAND2_X1 _07614_ ( .A1(_00662_ ), .A2(_00668_ ), .ZN(_00669_ ) );
NOR3_X1 _07615_ ( .A1(\u_idu.inst[5] ), .A2(\u_idu.inst[6] ), .A3(\u_idu.inst[4] ), .ZN(_00670_ ) );
AND2_X1 _07616_ ( .A1(_00665_ ), .A2(_00670_ ), .ZN(_00671_ ) );
OAI21_X1 _07617_ ( .A(\u_idu.imm_auipc_lui[13] ), .B1(\u_idu.imm_auipc_lui[12] ), .B2(\u_idu.imm_auipc_lui[14] ), .ZN(_00672_ ) );
AND2_X2 _07618_ ( .A1(_00671_ ), .A2(_00672_ ), .ZN(_00673_ ) );
INV_X1 _07619_ ( .A(_00673_ ), .ZN(_00674_ ) );
AND2_X1 _07620_ ( .A1(_00669_ ), .A2(_00674_ ), .ZN(_00675_ ) );
INV_X1 _07621_ ( .A(_00675_ ), .ZN(_00676_ ) );
INV_X1 _07622_ ( .A(\u_idu.imm_auipc_lui[13] ), .ZN(_00677_ ) );
OR3_X1 _07623_ ( .A1(_00645_ ), .A2(_00677_ ), .A3(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00678_ ) );
INV_X1 _07624_ ( .A(_00651_ ), .ZN(_00679_ ) );
OAI21_X1 _07625_ ( .A(_00678_ ), .B1(_00679_ ), .B2(_00647_ ), .ZN(_00680_ ) );
NOR3_X1 _07626_ ( .A1(_00677_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(\u_idu.imm_auipc_lui[12] ), .ZN(_00681_ ) );
AOI21_X1 _07627_ ( .A(_00681_ ), .B1(\u_idu.imm_auipc_lui[14] ), .B2(_00657_ ), .ZN(_00682_ ) );
INV_X1 _07628_ ( .A(_00682_ ), .ZN(_00683_ ) );
AND2_X2 _07629_ ( .A1(_00651_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00684_ ) );
NAND2_X1 _07630_ ( .A1(_00645_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00685_ ) );
NOR2_X1 _07631_ ( .A1(_00685_ ), .A2(\u_idu.imm_auipc_lui[13] ), .ZN(_00686_ ) );
BUF_X2 _07632_ ( .A(_00686_ ), .Z(_00687_ ) );
NOR4_X1 _07633_ ( .A1(_00680_ ), .A2(_00683_ ), .A3(_00684_ ), .A4(_00687_ ), .ZN(_00688_ ) );
INV_X1 _07634_ ( .A(\u_idu.inst[4] ), .ZN(_00689_ ) );
NAND2_X1 _07635_ ( .A1(_00689_ ), .A2(\u_idu.inst[5] ), .ZN(_00690_ ) );
NOR2_X1 _07636_ ( .A1(_00690_ ), .A2(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ), .ZN(_00691_ ) );
AND2_X2 _07637_ ( .A1(_00665_ ), .A2(_00691_ ), .ZN(_00692_ ) );
INV_X1 _07638_ ( .A(_00692_ ), .ZN(_00693_ ) );
NOR2_X1 _07639_ ( .A1(_00688_ ), .A2(_00693_ ), .ZN(_00694_ ) );
AND3_X1 _07640_ ( .A1(_00663_ ), .A2(\u_idu.inst[3] ), .A3(\u_idu.inst[2] ), .ZN(_00695_ ) );
AND2_X1 _07641_ ( .A1(_00695_ ), .A2(_00670_ ), .ZN(_00696_ ) );
INV_X1 _07642_ ( .A(_00696_ ), .ZN(_00697_ ) );
NOR2_X1 _07643_ ( .A1(_00697_ ), .A2(_00684_ ), .ZN(_00698_ ) );
NOR2_X1 _07644_ ( .A1(_00666_ ), .A2(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ), .ZN(_00699_ ) );
AND2_X2 _07645_ ( .A1(_00665_ ), .A2(_00699_ ), .ZN(_00700_ ) );
INV_X1 _07646_ ( .A(_00700_ ), .ZN(_00701_ ) );
NOR2_X1 _07647_ ( .A1(_00677_ ), .A2(\u_idu.imm_auipc_lui[12] ), .ZN(_00702_ ) );
AND2_X2 _07648_ ( .A1(_00702_ ), .A2(_00647_ ), .ZN(_00703_ ) );
NOR2_X1 _07649_ ( .A1(_00684_ ), .A2(_00703_ ), .ZN(_00704_ ) );
NOR2_X1 _07650_ ( .A1(_00701_ ), .A2(_00704_ ), .ZN(_00705_ ) );
NOR2_X1 _07651_ ( .A1(\u_idu.imm_auipc_lui[25] ), .A2(\u_idu.imm_auipc_lui[24] ), .ZN(_00706_ ) );
INV_X1 _07652_ ( .A(\u_idu.imm_auipc_lui[27] ), .ZN(_00707_ ) );
AND2_X1 _07653_ ( .A1(_00706_ ), .A2(_00707_ ), .ZN(_00708_ ) );
NOR2_X1 _07654_ ( .A1(\u_idu.imm_auipc_lui[23] ), .A2(\u_idu.imm_auipc_lui[26] ), .ZN(_00709_ ) );
AND2_X1 _07655_ ( .A1(_00708_ ), .A2(_00709_ ), .ZN(_00710_ ) );
NOR2_X1 _07656_ ( .A1(\u_idu.imm_auipc_lui[22] ), .A2(fanout_net_23 ), .ZN(_00711_ ) );
AND2_X1 _07657_ ( .A1(_00711_ ), .A2(fanout_net_22 ), .ZN(_00712_ ) );
AND2_X1 _07658_ ( .A1(_00638_ ), .A2(_00641_ ), .ZN(_00713_ ) );
NAND3_X1 _07659_ ( .A1(_00710_ ), .A2(_00712_ ), .A3(_00713_ ), .ZN(_00714_ ) );
INV_X1 _07660_ ( .A(_00686_ ), .ZN(_00715_ ) );
NOR2_X1 _07661_ ( .A1(_00714_ ), .A2(_00715_ ), .ZN(_00716_ ) );
AOI21_X1 _07662_ ( .A(_00705_ ), .B1(_00716_ ), .B2(_00700_ ), .ZN(_00717_ ) );
NAND3_X1 _07663_ ( .A1(\u_idu.inst[2] ), .A2(\u_idu.inst[0] ), .A3(\u_idu.inst[1] ), .ZN(_00718_ ) );
NOR2_X1 _07664_ ( .A1(_00718_ ), .A2(\u_idu.inst[3] ), .ZN(_00719_ ) );
AND2_X1 _07665_ ( .A1(_00691_ ), .A2(_00719_ ), .ZN(_00720_ ) );
AND2_X1 _07666_ ( .A1(_00720_ ), .A2(_00687_ ), .ZN(_00721_ ) );
INV_X1 _07667_ ( .A(_00721_ ), .ZN(_00722_ ) );
BUF_X2 _07668_ ( .A(_00722_ ), .Z(_00723_ ) );
INV_X1 _07669_ ( .A(\u_idu.inst[6] ), .ZN(_00724_ ) );
AND3_X1 _07670_ ( .A1(_00663_ ), .A2(_00724_ ), .A3(_00664_ ), .ZN(_00725_ ) );
AND2_X2 _07671_ ( .A1(_00725_ ), .A2(_00689_ ), .ZN(_00726_ ) );
AND2_X2 _07672_ ( .A1(_00726_ ), .A2(\u_idu.inst[5] ), .ZN(_00727_ ) );
INV_X1 _07673_ ( .A(_00727_ ), .ZN(_00728_ ) );
NOR3_X1 _07674_ ( .A1(_00684_ ), .A2(_00703_ ), .A3(_00686_ ), .ZN(_00729_ ) );
OAI211_X1 _07675_ ( .A(_00717_ ), .B(_00723_ ), .C1(_00728_ ), .C2(_00729_ ), .ZN(_00730_ ) );
OR4_X1 _07676_ ( .A1(_00676_ ), .A2(_00694_ ), .A3(_00698_ ), .A4(_00730_ ), .ZN(_00731_ ) );
NOR3_X1 _07677_ ( .A1(_00689_ ), .A2(\u_idu.inst[5] ), .A3(\u_idu.inst[6] ), .ZN(_00732_ ) );
AND2_X1 _07678_ ( .A1(_00665_ ), .A2(_00732_ ), .ZN(_00733_ ) );
BUF_X2 _07679_ ( .A(_00733_ ), .Z(_00734_ ) );
NOR2_X1 _07680_ ( .A1(_00731_ ), .A2(_00734_ ), .ZN(_00735_ ) );
INV_X1 _07681_ ( .A(_00735_ ), .ZN(_00736_ ) );
NOR2_X1 _07682_ ( .A1(_00689_ ), .A2(\u_idu.inst[6] ), .ZN(_00737_ ) );
AND2_X2 _07683_ ( .A1(_00719_ ), .A2(_00737_ ), .ZN(_00738_ ) );
NOR2_X1 _07684_ ( .A1(_00733_ ), .A2(_00738_ ), .ZN(_00739_ ) );
INV_X1 _07685_ ( .A(_00729_ ), .ZN(_00740_ ) );
AND2_X1 _07686_ ( .A1(_00727_ ), .A2(_00740_ ), .ZN(_00741_ ) );
AND2_X1 _07687_ ( .A1(_00696_ ), .A2(_00684_ ), .ZN(_00742_ ) );
BUF_X4 _07688_ ( .A(_00721_ ), .Z(_00743_ ) );
NOR4_X1 _07689_ ( .A1(_00741_ ), .A2(_00742_ ), .A3(_00705_ ), .A4(_00743_ ), .ZN(_00744_ ) );
NAND4_X1 _07690_ ( .A1(_00736_ ), .A2(_00675_ ), .A3(_00739_ ), .A4(_00744_ ), .ZN(_00745_ ) );
AND2_X2 _07691_ ( .A1(_00695_ ), .A2(_00691_ ), .ZN(_00746_ ) );
NOR2_X1 _07692_ ( .A1(_00721_ ), .A2(_00746_ ), .ZN(_00747_ ) );
INV_X1 _07693_ ( .A(fanout_net_23 ), .ZN(_00748_ ) );
NOR2_X1 _07694_ ( .A1(_00748_ ), .A2(\u_idu.imm_auipc_lui[22] ), .ZN(_00749_ ) );
INV_X1 _07695_ ( .A(\u_idu.imm_auipc_lui[23] ), .ZN(_00750_ ) );
INV_X1 _07696_ ( .A(fanout_net_22 ), .ZN(_00751_ ) );
AND3_X1 _07697_ ( .A1(_00749_ ), .A2(_00750_ ), .A3(_00751_ ), .ZN(_00752_ ) );
AND2_X1 _07698_ ( .A1(_00639_ ), .A2(_00706_ ), .ZN(_00753_ ) );
AND2_X1 _07699_ ( .A1(\u_idu.imm_auipc_lui[28] ), .A2(\u_idu.imm_auipc_lui[29] ), .ZN(_00754_ ) );
AND2_X2 _07700_ ( .A1(_00754_ ), .A2(_00641_ ), .ZN(_00755_ ) );
NAND3_X1 _07701_ ( .A1(_00752_ ), .A2(_00753_ ), .A3(_00755_ ), .ZN(_00756_ ) );
NOR2_X1 _07702_ ( .A1(_00756_ ), .A2(_00715_ ), .ZN(_00757_ ) );
NAND2_X1 _07703_ ( .A1(_00757_ ), .A2(_00700_ ), .ZN(_00758_ ) );
AND2_X1 _07704_ ( .A1(_00747_ ), .A2(_00758_ ), .ZN(_00759_ ) );
AND2_X1 _07705_ ( .A1(_00745_ ), .A2(_00759_ ), .ZN(_00760_ ) );
INV_X1 _07706_ ( .A(_00742_ ), .ZN(_00761_ ) );
AND2_X1 _07707_ ( .A1(_00760_ ), .A2(_00761_ ), .ZN(_00762_ ) );
INV_X1 _07708_ ( .A(_00632_ ), .ZN(_00763_ ) );
INV_X1 _07709_ ( .A(\u_exu.eopt[12] ), .ZN(_00764_ ) );
OR4_X1 _07710_ ( .A1(\ea_mask[1] ), .A2(_00764_ ), .A3(\ea_mask[0] ), .A4(\u_exu.eopt[15] ), .ZN(_00765_ ) );
NOR3_X2 _07711_ ( .A1(_00763_ ), .A2(\u_exu.eopt[0] ), .A3(_00765_ ), .ZN(_00766_ ) );
NOR2_X1 _07712_ ( .A1(_00766_ ), .A2(\u_exu.jmpc_ok ), .ZN(_00767_ ) );
OAI21_X1 _07713_ ( .A(_00637_ ), .B1(_00762_ ), .B2(_00767_ ), .ZN(_00768_ ) );
INV_X1 _07714_ ( .A(idu_ready ), .ZN(_00769_ ) );
NOR2_X2 _07715_ ( .A1(_00769_ ), .A2(exe_valid ), .ZN(_00770_ ) );
BUF_X4 _07716_ ( .A(_00770_ ), .Z(_00771_ ) );
OR2_X1 _07717_ ( .A1(_00768_ ), .A2(_00771_ ), .ZN(_00000_ ) );
INV_X1 _07718_ ( .A(fanout_net_1 ), .ZN(_00772_ ) );
BUF_X2 _07719_ ( .A(_00772_ ), .Z(_00773_ ) );
CLKBUF_X2 _07720_ ( .A(_00773_ ), .Z(_00774_ ) );
AND2_X1 _07721_ ( .A1(_00774_ ), .A2(\ea_addr[31] ), .ZN(_00001_ ) );
AND2_X1 _07722_ ( .A1(_00774_ ), .A2(\ea_addr[30] ), .ZN(_00002_ ) );
AND2_X1 _07723_ ( .A1(_00774_ ), .A2(\ea_addr[21] ), .ZN(_00003_ ) );
AND2_X1 _07724_ ( .A1(_00774_ ), .A2(\ea_addr[20] ), .ZN(_00004_ ) );
AND2_X1 _07725_ ( .A1(_00774_ ), .A2(\ea_addr[19] ), .ZN(_00005_ ) );
AND2_X1 _07726_ ( .A1(_00774_ ), .A2(\ea_addr[18] ), .ZN(_00006_ ) );
AND2_X1 _07727_ ( .A1(_00774_ ), .A2(\ea_addr[17] ), .ZN(_00007_ ) );
CLKBUF_X2 _07728_ ( .A(_00773_ ), .Z(_00775_ ) );
AND2_X1 _07729_ ( .A1(_00775_ ), .A2(\ea_addr[16] ), .ZN(_00008_ ) );
AND2_X1 _07730_ ( .A1(_00775_ ), .A2(\ea_addr[15] ), .ZN(_00009_ ) );
AND2_X1 _07731_ ( .A1(_00775_ ), .A2(\ea_addr[14] ), .ZN(_00010_ ) );
AND2_X1 _07732_ ( .A1(_00775_ ), .A2(\ea_addr[13] ), .ZN(_00011_ ) );
AND2_X1 _07733_ ( .A1(_00775_ ), .A2(\ea_addr[12] ), .ZN(_00012_ ) );
AND2_X1 _07734_ ( .A1(_00775_ ), .A2(\ea_addr[29] ), .ZN(_00013_ ) );
AND2_X1 _07735_ ( .A1(_00775_ ), .A2(\ea_addr[11] ), .ZN(_00014_ ) );
AND2_X1 _07736_ ( .A1(_00775_ ), .A2(\ea_addr[10] ), .ZN(_00015_ ) );
AND2_X1 _07737_ ( .A1(_00775_ ), .A2(\ea_addr[9] ), .ZN(_00016_ ) );
AND2_X1 _07738_ ( .A1(_00775_ ), .A2(\ea_addr[8] ), .ZN(_00017_ ) );
CLKBUF_X2 _07739_ ( .A(_00773_ ), .Z(_00776_ ) );
AND2_X1 _07740_ ( .A1(_00776_ ), .A2(\ea_addr[7] ), .ZN(_00018_ ) );
AND2_X1 _07741_ ( .A1(_00776_ ), .A2(\ea_addr[6] ), .ZN(_00019_ ) );
AND2_X1 _07742_ ( .A1(_00776_ ), .A2(\ea_addr[5] ), .ZN(_00020_ ) );
AND2_X1 _07743_ ( .A1(_00776_ ), .A2(\ea_addr[4] ), .ZN(_00021_ ) );
AND2_X1 _07744_ ( .A1(_00776_ ), .A2(\ea_addr[3] ), .ZN(_00022_ ) );
AND2_X1 _07745_ ( .A1(_00776_ ), .A2(\ea_addr[2] ), .ZN(_00023_ ) );
AND2_X1 _07746_ ( .A1(_00776_ ), .A2(\ea_addr[28] ), .ZN(_00024_ ) );
AND2_X1 _07747_ ( .A1(_00776_ ), .A2(\ea_addr[1] ), .ZN(_00025_ ) );
AND2_X1 _07748_ ( .A1(_00776_ ), .A2(\ea_addr[0] ), .ZN(_00026_ ) );
AND2_X1 _07749_ ( .A1(_00776_ ), .A2(\ea_addr[27] ), .ZN(_00027_ ) );
CLKBUF_X2 _07750_ ( .A(_00773_ ), .Z(_00777_ ) );
AND2_X1 _07751_ ( .A1(_00777_ ), .A2(\ea_addr[26] ), .ZN(_00028_ ) );
AND2_X1 _07752_ ( .A1(_00777_ ), .A2(\ea_addr[25] ), .ZN(_00029_ ) );
AND2_X1 _07753_ ( .A1(_00777_ ), .A2(\ea_addr[24] ), .ZN(_00030_ ) );
AND2_X1 _07754_ ( .A1(_00777_ ), .A2(\ea_addr[23] ), .ZN(_00031_ ) );
AND2_X1 _07755_ ( .A1(_00777_ ), .A2(\ea_addr[22] ), .ZN(_00032_ ) );
NOR2_X1 _07756_ ( .A1(_00627_ ), .A2(fanout_net_1 ), .ZN(_00033_ ) );
NOR2_X1 _07757_ ( .A1(_00628_ ), .A2(fanout_net_1 ), .ZN(_00034_ ) );
AND2_X1 _07758_ ( .A1(_00777_ ), .A2(ea_rsign ), .ZN(_00035_ ) );
AND2_X1 _07759_ ( .A1(_00629_ ), .A2(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ), .ZN(_00778_ ) );
AND3_X1 _07760_ ( .A1(_00632_ ), .A2(\u_exu.eopt[12] ), .A3(_00778_ ), .ZN(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_AND__A_Y ) );
CLKBUF_X2 _07761_ ( .A(_00772_ ), .Z(_00779_ ) );
AND4_X1 _07762_ ( .A1(_00779_ ), .A2(_00632_ ), .A3(\u_exu.eopt[12] ), .A4(_00778_ ), .ZN(_00036_ ) );
AND2_X1 _07763_ ( .A1(_00777_ ), .A2(\ea_ard[3] ), .ZN(_00037_ ) );
AND2_X1 _07764_ ( .A1(_00777_ ), .A2(\ea_ard[2] ), .ZN(_00038_ ) );
AND2_X1 _07765_ ( .A1(_00777_ ), .A2(\ea_ard[1] ), .ZN(_00039_ ) );
AND2_X1 _07766_ ( .A1(_00777_ ), .A2(\ea_ard[0] ), .ZN(_00040_ ) );
CLKBUF_X2 _07767_ ( .A(_00773_ ), .Z(_00780_ ) );
AND2_X1 _07768_ ( .A1(_00780_ ), .A2(\ea_wdata[31] ), .ZN(_00041_ ) );
AND2_X1 _07769_ ( .A1(_00780_ ), .A2(\ea_wdata[30] ), .ZN(_00042_ ) );
AND2_X1 _07770_ ( .A1(_00780_ ), .A2(\ea_wdata[21] ), .ZN(_00043_ ) );
AND2_X1 _07771_ ( .A1(_00780_ ), .A2(\ea_wdata[20] ), .ZN(_00044_ ) );
AND2_X1 _07772_ ( .A1(_00780_ ), .A2(\ea_wdata[19] ), .ZN(_00045_ ) );
AND2_X1 _07773_ ( .A1(_00780_ ), .A2(\ea_wdata[18] ), .ZN(_00046_ ) );
AND2_X1 _07774_ ( .A1(_00780_ ), .A2(\ea_wdata[17] ), .ZN(_00047_ ) );
AND2_X1 _07775_ ( .A1(_00780_ ), .A2(\ea_wdata[16] ), .ZN(_00048_ ) );
AND2_X1 _07776_ ( .A1(_00780_ ), .A2(\ea_wdata[15] ), .ZN(_00049_ ) );
AND2_X1 _07777_ ( .A1(_00780_ ), .A2(\ea_wdata[14] ), .ZN(_00050_ ) );
CLKBUF_X2 _07778_ ( .A(_00773_ ), .Z(_00781_ ) );
AND2_X1 _07779_ ( .A1(_00781_ ), .A2(\ea_wdata[13] ), .ZN(_00051_ ) );
AND2_X1 _07780_ ( .A1(_00781_ ), .A2(\ea_wdata[12] ), .ZN(_00052_ ) );
AND2_X1 _07781_ ( .A1(_00781_ ), .A2(\ea_wdata[29] ), .ZN(_00053_ ) );
AND2_X1 _07782_ ( .A1(_00781_ ), .A2(\ea_wdata[11] ), .ZN(_00054_ ) );
AND2_X1 _07783_ ( .A1(_00781_ ), .A2(\ea_wdata[10] ), .ZN(_00055_ ) );
AND2_X1 _07784_ ( .A1(_00781_ ), .A2(\ea_wdata[9] ), .ZN(_00056_ ) );
AND2_X1 _07785_ ( .A1(_00781_ ), .A2(\ea_wdata[8] ), .ZN(_00057_ ) );
AND2_X1 _07786_ ( .A1(_00781_ ), .A2(\ea_wdata[7] ), .ZN(_00058_ ) );
AND2_X1 _07787_ ( .A1(_00781_ ), .A2(\ea_wdata[6] ), .ZN(_00059_ ) );
AND2_X1 _07788_ ( .A1(_00781_ ), .A2(\ea_wdata[5] ), .ZN(_00060_ ) );
CLKBUF_X2 _07789_ ( .A(_00773_ ), .Z(_00782_ ) );
AND2_X1 _07790_ ( .A1(_00782_ ), .A2(\ea_wdata[4] ), .ZN(_00061_ ) );
AND2_X1 _07791_ ( .A1(_00782_ ), .A2(\ea_wdata[3] ), .ZN(_00062_ ) );
AND2_X1 _07792_ ( .A1(_00782_ ), .A2(\ea_wdata[2] ), .ZN(_00063_ ) );
AND2_X1 _07793_ ( .A1(_00782_ ), .A2(\ea_wdata[28] ), .ZN(_00064_ ) );
AND2_X1 _07794_ ( .A1(_00782_ ), .A2(\ea_wdata[1] ), .ZN(_00065_ ) );
AND2_X1 _07795_ ( .A1(_00782_ ), .A2(\ea_wdata[0] ), .ZN(_00066_ ) );
AND2_X1 _07796_ ( .A1(_00782_ ), .A2(\ea_wdata[27] ), .ZN(_00067_ ) );
AND2_X1 _07797_ ( .A1(_00782_ ), .A2(\ea_wdata[26] ), .ZN(_00068_ ) );
AND2_X1 _07798_ ( .A1(_00782_ ), .A2(\ea_wdata[25] ), .ZN(_00069_ ) );
AND2_X1 _07799_ ( .A1(_00782_ ), .A2(\ea_wdata[24] ), .ZN(_00070_ ) );
CLKBUF_X2 _07800_ ( .A(_00773_ ), .Z(_00783_ ) );
AND2_X1 _07801_ ( .A1(_00783_ ), .A2(\ea_wdata[23] ), .ZN(_00071_ ) );
AND2_X1 _07802_ ( .A1(_00783_ ), .A2(\ea_wdata[22] ), .ZN(_00072_ ) );
AND3_X1 _07803_ ( .A1(_00632_ ), .A2(_00783_ ), .A3(_00778_ ), .ZN(_00073_ ) );
AND3_X1 _07804_ ( .A1(_00632_ ), .A2(_00764_ ), .A3(_00778_ ), .ZN(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND4_X1 _07805_ ( .A1(_00779_ ), .A2(_00632_ ), .A3(_00764_ ), .A4(_00778_ ), .ZN(_00074_ ) );
INV_X1 _07806_ ( .A(fanout_net_5 ), .ZN(_00784_ ) );
CLKBUF_X2 _07807_ ( .A(_00784_ ), .Z(_00785_ ) );
CLKBUF_X2 _07808_ ( .A(_00785_ ), .Z(_00786_ ) );
CLKBUF_X2 _07809_ ( .A(_00786_ ), .Z(_00787_ ) );
OR2_X1 _07810_ ( .A1(_00787_ ), .A2(\ea_pc[31] ), .ZN(_00788_ ) );
OR2_X1 _07811_ ( .A1(\ea_addr[31] ), .A2(fanout_net_5 ), .ZN(_00789_ ) );
AND3_X1 _07812_ ( .A1(_00788_ ), .A2(_00783_ ), .A3(_00789_ ), .ZN(_00075_ ) );
OR2_X1 _07813_ ( .A1(_00786_ ), .A2(\ea_pc[30] ), .ZN(_00790_ ) );
OR2_X1 _07814_ ( .A1(\ea_addr[30] ), .A2(fanout_net_5 ), .ZN(_00791_ ) );
AND3_X1 _07815_ ( .A1(_00790_ ), .A2(_00783_ ), .A3(_00791_ ), .ZN(_00076_ ) );
NAND2_X1 _07816_ ( .A1(_00787_ ), .A2(\ea_addr[21] ), .ZN(_00792_ ) );
NAND2_X1 _07817_ ( .A1(fanout_net_5 ), .A2(\ea_pc[21] ), .ZN(_00793_ ) );
AOI21_X1 _07818_ ( .A(fanout_net_1 ), .B1(_00792_ ), .B2(_00793_ ), .ZN(_00077_ ) );
OR2_X1 _07819_ ( .A1(_00786_ ), .A2(\ea_pc[20] ), .ZN(_00794_ ) );
OR2_X1 _07820_ ( .A1(\ea_addr[20] ), .A2(fanout_net_5 ), .ZN(_00795_ ) );
AND3_X1 _07821_ ( .A1(_00794_ ), .A2(_00783_ ), .A3(_00795_ ), .ZN(_00078_ ) );
BUF_X2 _07822_ ( .A(_00786_ ), .Z(_00796_ ) );
BUF_X2 _07823_ ( .A(_00796_ ), .Z(_00797_ ) );
OR2_X1 _07824_ ( .A1(_00797_ ), .A2(\ea_pc[19] ), .ZN(_00798_ ) );
OR2_X1 _07825_ ( .A1(\ea_addr[19] ), .A2(fanout_net_5 ), .ZN(_00799_ ) );
AND3_X1 _07826_ ( .A1(_00798_ ), .A2(_00783_ ), .A3(_00799_ ), .ZN(_00079_ ) );
OR2_X1 _07827_ ( .A1(_00797_ ), .A2(\ea_pc[18] ), .ZN(_00800_ ) );
OR2_X1 _07828_ ( .A1(\ea_addr[18] ), .A2(fanout_net_5 ), .ZN(_00801_ ) );
AND3_X1 _07829_ ( .A1(_00800_ ), .A2(_00783_ ), .A3(_00801_ ), .ZN(_00080_ ) );
OR2_X1 _07830_ ( .A1(_00796_ ), .A2(\ea_pc[17] ), .ZN(_00802_ ) );
OR2_X1 _07831_ ( .A1(\ea_addr[17] ), .A2(fanout_net_5 ), .ZN(_00803_ ) );
AND3_X1 _07832_ ( .A1(_00802_ ), .A2(_00783_ ), .A3(_00803_ ), .ZN(_00081_ ) );
OR2_X1 _07833_ ( .A1(_00797_ ), .A2(\ea_pc[16] ), .ZN(_00804_ ) );
OR2_X1 _07834_ ( .A1(\ea_addr[16] ), .A2(fanout_net_5 ), .ZN(_00805_ ) );
AND3_X1 _07835_ ( .A1(_00804_ ), .A2(_00783_ ), .A3(_00805_ ), .ZN(_00082_ ) );
OR2_X1 _07836_ ( .A1(_00797_ ), .A2(\ea_pc[15] ), .ZN(_00806_ ) );
CLKBUF_X2 _07837_ ( .A(_00773_ ), .Z(_00807_ ) );
OR2_X1 _07838_ ( .A1(\ea_addr[15] ), .A2(fanout_net_5 ), .ZN(_00808_ ) );
AND3_X1 _07839_ ( .A1(_00806_ ), .A2(_00807_ ), .A3(_00808_ ), .ZN(_00083_ ) );
OR2_X1 _07840_ ( .A1(_00797_ ), .A2(\ea_pc[14] ), .ZN(_00809_ ) );
OR2_X1 _07841_ ( .A1(\ea_addr[14] ), .A2(fanout_net_5 ), .ZN(_00810_ ) );
AND3_X1 _07842_ ( .A1(_00809_ ), .A2(_00807_ ), .A3(_00810_ ), .ZN(_00084_ ) );
OR2_X1 _07843_ ( .A1(_00796_ ), .A2(\ea_pc[13] ), .ZN(_00811_ ) );
OR2_X1 _07844_ ( .A1(\ea_addr[13] ), .A2(fanout_net_5 ), .ZN(_00812_ ) );
AND3_X1 _07845_ ( .A1(_00811_ ), .A2(_00807_ ), .A3(_00812_ ), .ZN(_00085_ ) );
OR2_X1 _07846_ ( .A1(_00796_ ), .A2(\ea_pc[10] ), .ZN(_00813_ ) );
OR2_X1 _07847_ ( .A1(\ea_addr[10] ), .A2(fanout_net_5 ), .ZN(_00814_ ) );
AND3_X1 _07848_ ( .A1(_00813_ ), .A2(_00807_ ), .A3(_00814_ ), .ZN(_00086_ ) );
OR2_X1 _07849_ ( .A1(_00787_ ), .A2(\ea_pc[29] ), .ZN(_00815_ ) );
OR2_X1 _07850_ ( .A1(\ea_addr[29] ), .A2(fanout_net_5 ), .ZN(_00816_ ) );
AND3_X1 _07851_ ( .A1(_00815_ ), .A2(_00807_ ), .A3(_00816_ ), .ZN(_00087_ ) );
OR2_X1 _07852_ ( .A1(_00786_ ), .A2(\ea_pc[9] ), .ZN(_00817_ ) );
OR2_X1 _07853_ ( .A1(\ea_addr[9] ), .A2(fanout_net_5 ), .ZN(_00818_ ) );
AND3_X1 _07854_ ( .A1(_00817_ ), .A2(_00807_ ), .A3(_00818_ ), .ZN(_00088_ ) );
OR2_X1 _07855_ ( .A1(_00787_ ), .A2(\ea_pc[8] ), .ZN(_00819_ ) );
OR2_X1 _07856_ ( .A1(\ea_addr[8] ), .A2(fanout_net_5 ), .ZN(_00820_ ) );
AND3_X1 _07857_ ( .A1(_00819_ ), .A2(_00807_ ), .A3(_00820_ ), .ZN(_00089_ ) );
OR2_X1 _07858_ ( .A1(_00796_ ), .A2(\ea_pc[7] ), .ZN(_00821_ ) );
OR2_X1 _07859_ ( .A1(\ea_addr[7] ), .A2(fanout_net_5 ), .ZN(_00822_ ) );
AND3_X1 _07860_ ( .A1(_00821_ ), .A2(_00807_ ), .A3(_00822_ ), .ZN(_00090_ ) );
NAND2_X1 _07861_ ( .A1(_00787_ ), .A2(\ea_addr[6] ), .ZN(_00823_ ) );
NAND2_X1 _07862_ ( .A1(fanout_net_5 ), .A2(\ea_pc[6] ), .ZN(_00824_ ) );
AOI21_X1 _07863_ ( .A(fanout_net_1 ), .B1(_00823_ ), .B2(_00824_ ), .ZN(_00091_ ) );
NAND2_X1 _07864_ ( .A1(_00787_ ), .A2(\ea_addr[5] ), .ZN(_00825_ ) );
NAND2_X1 _07865_ ( .A1(fanout_net_5 ), .A2(\ea_pc[5] ), .ZN(_00826_ ) );
AOI21_X1 _07866_ ( .A(fanout_net_1 ), .B1(_00825_ ), .B2(_00826_ ), .ZN(_00092_ ) );
OR2_X1 _07867_ ( .A1(_00796_ ), .A2(\ea_pc[4] ), .ZN(_00827_ ) );
OR2_X1 _07868_ ( .A1(\ea_addr[4] ), .A2(fanout_net_5 ), .ZN(_00828_ ) );
AND3_X1 _07869_ ( .A1(_00827_ ), .A2(_00807_ ), .A3(_00828_ ), .ZN(_00093_ ) );
NAND2_X1 _07870_ ( .A1(_00796_ ), .A2(\ea_addr[3] ), .ZN(_00829_ ) );
NAND2_X1 _07871_ ( .A1(fanout_net_5 ), .A2(\ea_pc[3] ), .ZN(_00830_ ) );
AOI21_X1 _07872_ ( .A(fanout_net_1 ), .B1(_00829_ ), .B2(_00830_ ), .ZN(_00094_ ) );
NAND2_X1 _07873_ ( .A1(_00796_ ), .A2(\ea_addr[2] ), .ZN(_00831_ ) );
NAND2_X1 _07874_ ( .A1(fanout_net_5 ), .A2(\ea_pc[2] ), .ZN(_00832_ ) );
AOI21_X1 _07875_ ( .A(fanout_net_1 ), .B1(_00831_ ), .B2(_00832_ ), .ZN(_00095_ ) );
NAND2_X1 _07876_ ( .A1(_00797_ ), .A2(\ea_addr[1] ), .ZN(_00833_ ) );
NAND2_X1 _07877_ ( .A1(fanout_net_5 ), .A2(\ea_pc[1] ), .ZN(_00834_ ) );
AOI21_X1 _07878_ ( .A(fanout_net_1 ), .B1(_00833_ ), .B2(_00834_ ), .ZN(_00096_ ) );
NAND2_X1 _07879_ ( .A1(_00797_ ), .A2(\ea_addr[0] ), .ZN(_00835_ ) );
NAND2_X1 _07880_ ( .A1(fanout_net_5 ), .A2(\ea_pc[0] ), .ZN(_00836_ ) );
AOI21_X1 _07881_ ( .A(fanout_net_1 ), .B1(_00835_ ), .B2(_00836_ ), .ZN(_00097_ ) );
OR2_X1 _07882_ ( .A1(_00786_ ), .A2(\ea_pc[28] ), .ZN(_00837_ ) );
OR2_X1 _07883_ ( .A1(\ea_addr[28] ), .A2(fanout_net_5 ), .ZN(_00838_ ) );
AND3_X1 _07884_ ( .A1(_00837_ ), .A2(_00807_ ), .A3(_00838_ ), .ZN(_00098_ ) );
OR2_X1 _07885_ ( .A1(_00787_ ), .A2(\ea_pc[27] ), .ZN(_00839_ ) );
CLKBUF_X2 _07886_ ( .A(_00773_ ), .Z(_00840_ ) );
OR2_X1 _07887_ ( .A1(\ea_addr[27] ), .A2(fanout_net_5 ), .ZN(_00841_ ) );
AND3_X1 _07888_ ( .A1(_00839_ ), .A2(_00840_ ), .A3(_00841_ ), .ZN(_00099_ ) );
OR2_X1 _07889_ ( .A1(_00787_ ), .A2(\ea_pc[26] ), .ZN(_00842_ ) );
OR2_X1 _07890_ ( .A1(\ea_addr[26] ), .A2(fanout_net_5 ), .ZN(_00843_ ) );
AND3_X1 _07891_ ( .A1(_00842_ ), .A2(_00840_ ), .A3(_00843_ ), .ZN(_00100_ ) );
OR2_X1 _07892_ ( .A1(_00786_ ), .A2(\ea_pc[25] ), .ZN(_00844_ ) );
OR2_X1 _07893_ ( .A1(\ea_addr[25] ), .A2(fanout_net_5 ), .ZN(_00845_ ) );
AND3_X1 _07894_ ( .A1(_00844_ ), .A2(_00840_ ), .A3(_00845_ ), .ZN(_00101_ ) );
NAND2_X1 _07895_ ( .A1(_00787_ ), .A2(\ea_addr[24] ), .ZN(_00846_ ) );
NAND2_X1 _07896_ ( .A1(ea_err ), .A2(\ea_pc[24] ), .ZN(_00847_ ) );
AOI21_X1 _07897_ ( .A(fanout_net_1 ), .B1(_00846_ ), .B2(_00847_ ), .ZN(_00102_ ) );
OR2_X1 _07898_ ( .A1(_00786_ ), .A2(\ea_pc[23] ), .ZN(_00848_ ) );
OR2_X1 _07899_ ( .A1(\ea_addr[23] ), .A2(ea_err ), .ZN(_00849_ ) );
AND3_X1 _07900_ ( .A1(_00848_ ), .A2(_00840_ ), .A3(_00849_ ), .ZN(_00103_ ) );
OR2_X1 _07901_ ( .A1(_00787_ ), .A2(\ea_pc[22] ), .ZN(_00850_ ) );
OR2_X1 _07902_ ( .A1(\ea_addr[22] ), .A2(ea_err ), .ZN(_00851_ ) );
AND3_X1 _07903_ ( .A1(_00850_ ), .A2(_00840_ ), .A3(_00851_ ), .ZN(_00104_ ) );
NAND2_X1 _07904_ ( .A1(_00796_ ), .A2(\ea_addr[12] ), .ZN(_00852_ ) );
NAND2_X1 _07905_ ( .A1(ea_err ), .A2(\ea_pc[12] ), .ZN(_00853_ ) );
NAND3_X1 _07906_ ( .A1(_00852_ ), .A2(_00774_ ), .A3(_00853_ ), .ZN(_00105_ ) );
NAND2_X1 _07907_ ( .A1(_00797_ ), .A2(\ea_addr[11] ), .ZN(_00854_ ) );
NAND2_X1 _07908_ ( .A1(ea_err ), .A2(\ea_pc[11] ), .ZN(_00855_ ) );
NAND3_X1 _07909_ ( .A1(_00854_ ), .A2(_00774_ ), .A3(_00855_ ), .ZN(_00106_ ) );
AOI21_X1 _07910_ ( .A(fanout_net_1 ), .B1(_00852_ ), .B2(_00853_ ), .ZN(_00107_ ) );
AOI21_X1 _07911_ ( .A(fanout_net_1 ), .B1(_00854_ ), .B2(_00855_ ), .ZN(_00108_ ) );
BUF_X8 _07912_ ( .A(_00766_ ), .Z(_00856_ ) );
BUF_X4 _07913_ ( .A(_00856_ ), .Z(_00857_ ) );
BUF_X4 _07914_ ( .A(_00634_ ), .Z(_00858_ ) );
BUF_X4 _07915_ ( .A(_00858_ ), .Z(_00859_ ) );
BUF_X4 _07916_ ( .A(_00859_ ), .Z(_00860_ ) );
NOR4_X1 _07917_ ( .A1(_00857_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00653_ ), .ZN(_00110_ ) );
BUF_X4 _07918_ ( .A(_00856_ ), .Z(_00861_ ) );
INV_X1 _07919_ ( .A(\u_idu.imm_auipc_lui[30] ), .ZN(_00862_ ) );
NOR4_X1 _07920_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00862_ ), .ZN(_00111_ ) );
NOR2_X1 _07921_ ( .A1(_00766_ ), .A2(fanout_net_1 ), .ZN(_00863_ ) );
BUF_X2 _07922_ ( .A(_00863_ ), .Z(_00864_ ) );
CLKBUF_X2 _07923_ ( .A(_00864_ ), .Z(_00865_ ) );
CLKBUF_X2 _07924_ ( .A(_00637_ ), .Z(_00866_ ) );
AND4_X1 _07925_ ( .A1(_00750_ ), .A2(_00755_ ), .A3(_00753_ ), .A4(_00749_ ), .ZN(_00867_ ) );
AND2_X1 _07926_ ( .A1(_00686_ ), .A2(\u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ), .ZN(_00868_ ) );
NAND2_X1 _07927_ ( .A1(_00867_ ), .A2(_00868_ ), .ZN(_00869_ ) );
NAND4_X1 _07928_ ( .A1(_00710_ ), .A2(_00686_ ), .A3(_00712_ ), .A4(_00713_ ), .ZN(_00870_ ) );
AND2_X1 _07929_ ( .A1(_00869_ ), .A2(_00870_ ), .ZN(_00871_ ) );
AND2_X1 _07930_ ( .A1(_00871_ ), .A2(fanout_net_23 ), .ZN(_00872_ ) );
AND3_X1 _07931_ ( .A1(_00865_ ), .A2(_00866_ ), .A3(_00872_ ), .ZN(_00112_ ) );
NOR2_X1 _07932_ ( .A1(_00858_ ), .A2(fanout_net_1 ), .ZN(_00873_ ) );
INV_X2 _07933_ ( .A(_00873_ ), .ZN(_00874_ ) );
BUF_X2 _07934_ ( .A(_00874_ ), .Z(flush_$_OR__Y_B ) );
BUF_X2 _07935_ ( .A(_00751_ ), .Z(_00875_ ) );
BUF_X4 _07936_ ( .A(_00875_ ), .Z(_00876_ ) );
BUF_X4 _07937_ ( .A(_00876_ ), .Z(_00877_ ) );
BUF_X4 _07938_ ( .A(_00877_ ), .Z(_00878_ ) );
BUF_X4 _07939_ ( .A(_00766_ ), .Z(_00879_ ) );
INV_X1 _07940_ ( .A(\u_idu.imm_auipc_lui[26] ), .ZN(_00880_ ) );
NAND4_X1 _07941_ ( .A1(_00749_ ), .A2(_00750_ ), .A3(_00880_ ), .A4(_00706_ ), .ZN(_00881_ ) );
INV_X1 _07942_ ( .A(\u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ), .ZN(_00882_ ) );
NOR3_X1 _07943_ ( .A1(_00715_ ), .A2(_00881_ ), .A3(_00882_ ), .ZN(_00883_ ) );
AND3_X1 _07944_ ( .A1(_00754_ ), .A2(_00707_ ), .A3(_00641_ ), .ZN(_00884_ ) );
AND2_X1 _07945_ ( .A1(_00883_ ), .A2(_00884_ ), .ZN(_00885_ ) );
AND3_X1 _07946_ ( .A1(_00753_ ), .A2(_00712_ ), .A3(_00750_ ), .ZN(_00886_ ) );
AND3_X1 _07947_ ( .A1(_00886_ ), .A2(_00687_ ), .A3(_00713_ ), .ZN(_00887_ ) );
OR2_X1 _07948_ ( .A1(_00885_ ), .A2(_00887_ ), .ZN(_00888_ ) );
NOR4_X1 _07949_ ( .A1(flush_$_OR__Y_B ), .A2(_00878_ ), .A3(_00879_ ), .A4(_00888_ ), .ZN(_00113_ ) );
INV_X1 _07950_ ( .A(\u_idu.imm_auipc_lui[29] ), .ZN(_00889_ ) );
NOR4_X1 _07951_ ( .A1(flush_$_OR__Y_B ), .A2(_00889_ ), .A3(_00879_ ), .A4(_00888_ ), .ZN(_00114_ ) );
INV_X1 _07952_ ( .A(\u_idu.imm_auipc_lui[28] ), .ZN(_00890_ ) );
NOR4_X1 _07953_ ( .A1(flush_$_OR__Y_B ), .A2(_00890_ ), .A3(_00879_ ), .A4(_00888_ ), .ZN(_00115_ ) );
NOR4_X1 _07954_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00707_ ), .ZN(_00116_ ) );
NOR4_X1 _07955_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00880_ ), .ZN(_00117_ ) );
INV_X1 _07956_ ( .A(\u_idu.imm_auipc_lui[25] ), .ZN(_00891_ ) );
NOR4_X1 _07957_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00891_ ), .ZN(_00118_ ) );
INV_X1 _07958_ ( .A(\u_idu.imm_auipc_lui[24] ), .ZN(_00892_ ) );
NOR4_X1 _07959_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00892_ ), .ZN(_00119_ ) );
BUF_X2 _07960_ ( .A(_00750_ ), .Z(_00893_ ) );
NOR4_X1 _07961_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00893_ ), .ZN(_00120_ ) );
INV_X1 _07962_ ( .A(\u_idu.imm_auipc_lui[22] ), .ZN(_00894_ ) );
NOR4_X1 _07963_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_00894_ ), .ZN(_00121_ ) );
NOR2_X1 _07964_ ( .A1(_00874_ ), .A2(_00766_ ), .ZN(_00895_ ) );
INV_X2 _07965_ ( .A(_00895_ ), .ZN(_00896_ ) );
BUF_X4 _07966_ ( .A(_00896_ ), .Z(_00897_ ) );
BUF_X4 _07967_ ( .A(_00897_ ), .Z(_00898_ ) );
NOR3_X1 _07968_ ( .A1(_00668_ ), .A2(_00733_ ), .A3(_00720_ ), .ZN(_00899_ ) );
NOR2_X1 _07969_ ( .A1(_00726_ ), .A2(_00692_ ), .ZN(_00900_ ) );
AND2_X1 _07970_ ( .A1(_00899_ ), .A2(_00900_ ), .ZN(_00901_ ) );
OAI21_X2 _07971_ ( .A(_00901_ ), .B1(_00686_ ), .B2(_00701_ ), .ZN(_00902_ ) );
AND2_X1 _07972_ ( .A1(_00902_ ), .A2(fanout_net_21 ), .ZN(_00903_ ) );
BUF_X4 _07973_ ( .A(_00903_ ), .Z(_00904_ ) );
AOI21_X1 _07974_ ( .A(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ), .B1(_00899_ ), .B2(_00900_ ), .ZN(_00905_ ) );
AOI21_X1 _07975_ ( .A(_00701_ ), .B1(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ), .B2(_00715_ ), .ZN(_00906_ ) );
OR2_X2 _07976_ ( .A1(_00905_ ), .A2(_00906_ ), .ZN(_00907_ ) );
INV_X1 _07977_ ( .A(_00907_ ), .ZN(_00908_ ) );
NOR2_X2 _07978_ ( .A1(_00904_ ), .A2(_00908_ ), .ZN(_00909_ ) );
NAND2_X1 _07979_ ( .A1(_00901_ ), .A2(_00701_ ), .ZN(_00910_ ) );
OAI21_X1 _07980_ ( .A(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_B ), .B1(_00701_ ), .B2(_00715_ ), .ZN(_00911_ ) );
NAND2_X2 _07981_ ( .A1(_00910_ ), .A2(_00911_ ), .ZN(_00912_ ) );
INV_X1 _07982_ ( .A(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_1_B ), .ZN(_00913_ ) );
AND2_X1 _07983_ ( .A1(_00902_ ), .A2(_00913_ ), .ZN(_00914_ ) );
BUF_X4 _07984_ ( .A(_00914_ ), .Z(_00915_ ) );
NAND3_X1 _07985_ ( .A1(_00909_ ), .A2(_00912_ ), .A3(_00915_ ), .ZN(_00916_ ) );
AOI21_X1 _07986_ ( .A(_00668_ ), .B1(_00726_ ), .B2(\u_idu.inst[5] ), .ZN(_00917_ ) );
AND2_X1 _07987_ ( .A1(_00917_ ), .A2(_00693_ ), .ZN(_00918_ ) );
NOR2_X1 _07988_ ( .A1(_00918_ ), .A2(_00748_ ), .ZN(_00919_ ) );
AND2_X2 _07989_ ( .A1(_00919_ ), .A2(_00751_ ), .ZN(_00920_ ) );
NOR2_X1 _07990_ ( .A1(_00918_ ), .A2(_00894_ ), .ZN(_00921_ ) );
NAND3_X1 _07991_ ( .A1(_00920_ ), .A2(_00893_ ), .A3(_00921_ ), .ZN(_00922_ ) );
NAND2_X1 _07992_ ( .A1(_00916_ ), .A2(_00922_ ), .ZN(_00923_ ) );
NOR2_X1 _07993_ ( .A1(_00746_ ), .A2(_00671_ ), .ZN(_00924_ ) );
INV_X1 _07994_ ( .A(_00668_ ), .ZN(_00925_ ) );
NAND3_X1 _07995_ ( .A1(_00924_ ), .A2(_00925_ ), .A3(_00701_ ), .ZN(_00926_ ) );
INV_X1 _07996_ ( .A(_00733_ ), .ZN(_00927_ ) );
INV_X1 _07997_ ( .A(_00738_ ), .ZN(_00928_ ) );
INV_X1 _07998_ ( .A(_00720_ ), .ZN(_00929_ ) );
NAND3_X1 _07999_ ( .A1(_00927_ ), .A2(_00928_ ), .A3(_00929_ ), .ZN(_00930_ ) );
OAI21_X1 _08000_ ( .A(\u_idu.imm_branch[2] ), .B1(_00926_ ), .B2(_00930_ ), .ZN(_00931_ ) );
OR2_X1 _08001_ ( .A1(_00697_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00932_ ) );
AND2_X2 _08002_ ( .A1(_00931_ ), .A2(_00932_ ), .ZN(_00933_ ) );
INV_X1 _08003_ ( .A(_00933_ ), .ZN(_00934_ ) );
OAI21_X1 _08004_ ( .A(\u_idu.imm_branch[1] ), .B1(_00926_ ), .B2(_00930_ ), .ZN(_00935_ ) );
OR2_X1 _08005_ ( .A1(_00697_ ), .A2(de_ard_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00936_ ) );
AND2_X2 _08006_ ( .A1(_00935_ ), .A2(_00936_ ), .ZN(_00937_ ) );
INV_X1 _08007_ ( .A(_00937_ ), .ZN(_00938_ ) );
OAI21_X1 _08008_ ( .A(\u_idu.imm_branch[11] ), .B1(_00926_ ), .B2(_00930_ ), .ZN(_00939_ ) );
NAND3_X1 _08009_ ( .A1(_00695_ ), .A2(\u_idu.imm_auipc_lui[12] ), .A3(_00670_ ), .ZN(_00940_ ) );
AND2_X2 _08010_ ( .A1(_00939_ ), .A2(_00940_ ), .ZN(_00941_ ) );
NAND3_X1 _08011_ ( .A1(_00934_ ), .A2(_00938_ ), .A3(_00941_ ), .ZN(_00942_ ) );
NOR2_X1 _08012_ ( .A1(_00926_ ), .A2(_00930_ ), .ZN(_00943_ ) );
INV_X1 _08013_ ( .A(\u_idu.imm_branch[3] ), .ZN(_00944_ ) );
NOR2_X1 _08014_ ( .A1(_00943_ ), .A2(_00944_ ), .ZN(_00945_ ) );
BUF_X4 _08015_ ( .A(_00945_ ), .Z(_00946_ ) );
NOR2_X1 _08016_ ( .A1(_00942_ ), .A2(_00946_ ), .ZN(_00947_ ) );
OAI21_X1 _08017_ ( .A(\u_exu.rlock[6] ), .B1(_00923_ ), .B2(_00947_ ), .ZN(_00948_ ) );
AND2_X1 _08018_ ( .A1(_00904_ ), .A2(_00907_ ), .ZN(_00949_ ) );
BUF_X4 _08019_ ( .A(_00949_ ), .Z(_00950_ ) );
INV_X1 _08020_ ( .A(_00912_ ), .ZN(_00951_ ) );
INV_X1 _08021_ ( .A(_00914_ ), .ZN(_00952_ ) );
NAND3_X1 _08022_ ( .A1(_00950_ ), .A2(_00951_ ), .A3(_00952_ ), .ZN(_00953_ ) );
NOR2_X1 _08023_ ( .A1(_00918_ ), .A2(_00751_ ), .ZN(_00954_ ) );
BUF_X4 _08024_ ( .A(_00954_ ), .Z(_00955_ ) );
NAND3_X1 _08025_ ( .A1(_00955_ ), .A2(_00894_ ), .A3(fanout_net_23 ), .ZN(_00956_ ) );
OAI21_X1 _08026_ ( .A(_00953_ ), .B1(_00893_ ), .B2(_00956_ ), .ZN(_00957_ ) );
INV_X1 _08027_ ( .A(_00941_ ), .ZN(_00958_ ) );
NAND3_X1 _08028_ ( .A1(_00938_ ), .A2(_00958_ ), .A3(_00933_ ), .ZN(_00959_ ) );
INV_X2 _08029_ ( .A(_00945_ ), .ZN(_00960_ ) );
NOR2_X1 _08030_ ( .A1(_00959_ ), .A2(_00960_ ), .ZN(_00961_ ) );
OAI21_X1 _08031_ ( .A(\u_exu.rlock[11] ), .B1(_00957_ ), .B2(_00961_ ), .ZN(_00962_ ) );
NAND3_X1 _08032_ ( .A1(_00950_ ), .A2(_00951_ ), .A3(_00914_ ), .ZN(_00963_ ) );
NOR2_X1 _08033_ ( .A1(_00918_ ), .A2(_00893_ ), .ZN(_00964_ ) );
NAND4_X1 _08034_ ( .A1(_00964_ ), .A2(_00955_ ), .A3(\u_idu.imm_auipc_lui[22] ), .A4(fanout_net_23 ), .ZN(_00965_ ) );
NAND2_X1 _08035_ ( .A1(_00963_ ), .A2(_00965_ ), .ZN(_00966_ ) );
NAND3_X1 _08036_ ( .A1(_00934_ ), .A2(_00938_ ), .A3(_00958_ ), .ZN(_00967_ ) );
NOR2_X1 _08037_ ( .A1(_00967_ ), .A2(_00960_ ), .ZN(_00968_ ) );
OAI21_X1 _08038_ ( .A(\u_exu.rlock[15] ), .B1(_00966_ ), .B2(_00968_ ), .ZN(_00969_ ) );
NAND2_X1 _08039_ ( .A1(_00962_ ), .A2(_00969_ ), .ZN(_00970_ ) );
INV_X1 _08040_ ( .A(_00964_ ), .ZN(_00971_ ) );
INV_X1 _08041_ ( .A(_00921_ ), .ZN(_00972_ ) );
NAND3_X1 _08042_ ( .A1(_00920_ ), .A2(_00971_ ), .A3(_00972_ ), .ZN(_00973_ ) );
NAND3_X1 _08043_ ( .A1(_00938_ ), .A2(_00933_ ), .A3(_00941_ ), .ZN(_00974_ ) );
BUF_X4 _08044_ ( .A(_00952_ ), .Z(_00975_ ) );
INV_X1 _08045_ ( .A(_00904_ ), .ZN(_00976_ ) );
NAND3_X1 _08046_ ( .A1(_00975_ ), .A2(_00976_ ), .A3(_00907_ ), .ZN(_00977_ ) );
OAI221_X1 _08047_ ( .A(_00973_ ), .B1(_00946_ ), .B2(_00974_ ), .C1(_00977_ ), .C2(_00951_ ), .ZN(_00978_ ) );
NAND3_X1 _08048_ ( .A1(_00952_ ), .A2(_00976_ ), .A3(_00908_ ), .ZN(_00979_ ) );
INV_X1 _08049_ ( .A(_00919_ ), .ZN(_00980_ ) );
INV_X1 _08050_ ( .A(_00954_ ), .ZN(_00981_ ) );
NAND3_X1 _08051_ ( .A1(_00972_ ), .A2(_00980_ ), .A3(_00981_ ), .ZN(_00982_ ) );
OAI22_X1 _08052_ ( .A1(_00979_ ), .A2(_00951_ ), .B1(_00964_ ), .B2(_00982_ ), .ZN(_00983_ ) );
NAND3_X1 _08053_ ( .A1(_00933_ ), .A2(_00937_ ), .A3(_00941_ ), .ZN(_00984_ ) );
NOR2_X1 _08054_ ( .A1(_00984_ ), .A2(_00945_ ), .ZN(_00985_ ) );
OR2_X1 _08055_ ( .A1(_00983_ ), .A2(_00985_ ), .ZN(_00986_ ) );
AOI221_X4 _08056_ ( .A(_00970_ ), .B1(\u_exu.rlock[2] ), .B2(_00978_ ), .C1(\u_exu.rlock[0] ), .C2(_00986_ ), .ZN(_00987_ ) );
NOR2_X1 _08057_ ( .A1(_00919_ ), .A2(_00955_ ), .ZN(_00988_ ) );
NAND3_X1 _08058_ ( .A1(_00988_ ), .A2(_00964_ ), .A3(_00921_ ), .ZN(_00989_ ) );
NAND3_X1 _08059_ ( .A1(_00976_ ), .A2(_00914_ ), .A3(_00908_ ), .ZN(_00990_ ) );
OAI21_X1 _08060_ ( .A(_00989_ ), .B1(_00990_ ), .B2(_00912_ ), .ZN(_00991_ ) );
NAND3_X1 _08061_ ( .A1(_00934_ ), .A2(_00937_ ), .A3(_00941_ ), .ZN(_00992_ ) );
NOR2_X1 _08062_ ( .A1(_00992_ ), .A2(_00960_ ), .ZN(_00993_ ) );
OAI21_X1 _08063_ ( .A(\u_exu.rlock[12] ), .B1(_00991_ ), .B2(_00993_ ), .ZN(_00994_ ) );
AND2_X1 _08064_ ( .A1(_00954_ ), .A2(_00748_ ), .ZN(_00995_ ) );
BUF_X4 _08065_ ( .A(_00995_ ), .Z(_00996_ ) );
NAND3_X1 _08066_ ( .A1(_00996_ ), .A2(\u_idu.imm_auipc_lui[22] ), .A3(_00971_ ), .ZN(_00997_ ) );
NAND3_X1 _08067_ ( .A1(_00915_ ), .A2(_00904_ ), .A3(_00908_ ), .ZN(_00998_ ) );
OAI21_X1 _08068_ ( .A(_00997_ ), .B1(_00998_ ), .B2(_00951_ ), .ZN(_00999_ ) );
NAND3_X1 _08069_ ( .A1(_00934_ ), .A2(_00958_ ), .A3(_00937_ ), .ZN(_01000_ ) );
NOR2_X1 _08070_ ( .A1(_01000_ ), .A2(_00946_ ), .ZN(_01001_ ) );
OAI21_X1 _08071_ ( .A(\u_exu.rlock[5] ), .B1(_00999_ ), .B2(_01001_ ), .ZN(_01002_ ) );
AND2_X1 _08072_ ( .A1(_00994_ ), .A2(_01002_ ), .ZN(_01003_ ) );
AND2_X1 _08073_ ( .A1(_00904_ ), .A2(_00908_ ), .ZN(_01004_ ) );
BUF_X4 _08074_ ( .A(_01004_ ), .Z(_01005_ ) );
NAND3_X1 _08075_ ( .A1(_01005_ ), .A2(_00912_ ), .A3(_00975_ ), .ZN(_01006_ ) );
NAND3_X1 _08076_ ( .A1(_00958_ ), .A2(_00933_ ), .A3(_00937_ ), .ZN(_01007_ ) );
OAI21_X1 _08077_ ( .A(_01006_ ), .B1(_00946_ ), .B2(_01007_ ), .ZN(_01008_ ) );
AND4_X1 _08078_ ( .A1(_00971_ ), .A2(_00972_ ), .A3(_00980_ ), .A4(_00955_ ), .ZN(_01009_ ) );
OAI21_X1 _08079_ ( .A(\u_exu.rlock[1] ), .B1(_01008_ ), .B2(_01009_ ), .ZN(_01010_ ) );
NAND3_X1 _08080_ ( .A1(_00950_ ), .A2(_00912_ ), .A3(_00975_ ), .ZN(_01011_ ) );
OAI21_X1 _08081_ ( .A(_01011_ ), .B1(\u_idu.imm_auipc_lui[23] ), .B2(_00956_ ), .ZN(_01012_ ) );
NOR2_X1 _08082_ ( .A1(_00959_ ), .A2(_00946_ ), .ZN(_01013_ ) );
OAI21_X1 _08083_ ( .A(\u_exu.rlock[3] ), .B1(_01012_ ), .B2(_01013_ ), .ZN(_01014_ ) );
NAND3_X1 _08084_ ( .A1(_00996_ ), .A2(\u_idu.imm_auipc_lui[22] ), .A3(_00964_ ), .ZN(_01015_ ) );
OAI21_X1 _08085_ ( .A(_01015_ ), .B1(_00998_ ), .B2(_00912_ ), .ZN(_01016_ ) );
NOR2_X1 _08086_ ( .A1(_01000_ ), .A2(_00960_ ), .ZN(_01017_ ) );
OAI21_X1 _08087_ ( .A(\u_exu.rlock[13] ), .B1(_01016_ ), .B2(_01017_ ), .ZN(_01018_ ) );
AND3_X1 _08088_ ( .A1(_00909_ ), .A2(_00951_ ), .A3(_00915_ ), .ZN(_01019_ ) );
NAND3_X1 _08089_ ( .A1(_00920_ ), .A2(\u_idu.imm_auipc_lui[23] ), .A3(_00921_ ), .ZN(_01020_ ) );
OAI21_X1 _08090_ ( .A(_01020_ ), .B1(_00942_ ), .B2(_00960_ ), .ZN(_01021_ ) );
OAI21_X1 _08091_ ( .A(\u_exu.rlock[14] ), .B1(_01019_ ), .B2(_01021_ ), .ZN(_01022_ ) );
AND4_X1 _08092_ ( .A1(_01010_ ), .A2(_01014_ ), .A3(_01018_ ), .A4(_01022_ ), .ZN(_01023_ ) );
AND4_X1 _08093_ ( .A1(_00948_ ), .A2(_00987_ ), .A3(_01003_ ), .A4(_01023_ ), .ZN(_01024_ ) );
INV_X1 _08094_ ( .A(\u_exu.exe_start ), .ZN(_01025_ ) );
NAND3_X1 _08095_ ( .A1(_01005_ ), .A2(_00951_ ), .A3(_00975_ ), .ZN(_01026_ ) );
NAND2_X1 _08096_ ( .A1(_00964_ ), .A2(_00712_ ), .ZN(_01027_ ) );
NAND2_X1 _08097_ ( .A1(_01026_ ), .A2(_01027_ ), .ZN(_01028_ ) );
NOR2_X1 _08098_ ( .A1(_01007_ ), .A2(_00960_ ), .ZN(_01029_ ) );
OAI21_X1 _08099_ ( .A(\u_exu.rlock[9] ), .B1(_01028_ ), .B2(_01029_ ), .ZN(_01030_ ) );
NAND3_X1 _08100_ ( .A1(_00950_ ), .A2(_00912_ ), .A3(_00915_ ), .ZN(_01031_ ) );
NAND4_X1 _08101_ ( .A1(_00971_ ), .A2(\u_idu.imm_auipc_lui[22] ), .A3(fanout_net_23 ), .A4(_00955_ ), .ZN(_01032_ ) );
NAND2_X1 _08102_ ( .A1(_01031_ ), .A2(_01032_ ), .ZN(_01033_ ) );
NOR2_X1 _08103_ ( .A1(_00967_ ), .A2(_00946_ ), .ZN(_01034_ ) );
OAI21_X1 _08104_ ( .A(\u_exu.rlock[7] ), .B1(_01033_ ), .B2(_01034_ ), .ZN(_01035_ ) );
OAI22_X1 _08105_ ( .A1(_00979_ ), .A2(_00912_ ), .B1(_00971_ ), .B2(_00982_ ), .ZN(_01036_ ) );
NOR2_X1 _08106_ ( .A1(_00984_ ), .A2(_00960_ ), .ZN(_01037_ ) );
OAI21_X1 _08107_ ( .A(\u_exu.rlock[8] ), .B1(_01036_ ), .B2(_01037_ ), .ZN(_01038_ ) );
NAND3_X1 _08108_ ( .A1(_00988_ ), .A2(_00971_ ), .A3(_00921_ ), .ZN(_01039_ ) );
OAI21_X1 _08109_ ( .A(_01039_ ), .B1(_00990_ ), .B2(_00951_ ), .ZN(_01040_ ) );
NOR2_X1 _08110_ ( .A1(_00992_ ), .A2(_00946_ ), .ZN(_01041_ ) );
OAI21_X1 _08111_ ( .A(\u_exu.rlock[4] ), .B1(_01040_ ), .B2(_01041_ ), .ZN(_01042_ ) );
AND4_X1 _08112_ ( .A1(_01030_ ), .A2(_01035_ ), .A3(_01038_ ), .A4(_01042_ ), .ZN(_01043_ ) );
BUF_X2 _08113_ ( .A(_00964_ ), .Z(_01044_ ) );
NAND3_X1 _08114_ ( .A1(_00920_ ), .A2(_01044_ ), .A3(_00972_ ), .ZN(_01045_ ) );
CLKBUF_X2 _08115_ ( .A(_00912_ ), .Z(_01046_ ) );
OAI221_X1 _08116_ ( .A(_01045_ ), .B1(_00960_ ), .B2(_00974_ ), .C1(_00977_ ), .C2(_01046_ ), .ZN(_01047_ ) );
NAND2_X1 _08117_ ( .A1(_01047_ ), .A2(\u_exu.rlock[10] ), .ZN(_01048_ ) );
AND4_X1 _08118_ ( .A1(_01025_ ), .A2(_01043_ ), .A3(exe_valid ), .A4(_01048_ ), .ZN(_01049_ ) );
AND2_X1 _08119_ ( .A1(_01024_ ), .A2(_01049_ ), .ZN(_01050_ ) );
INV_X1 _08120_ ( .A(_01050_ ), .ZN(_01051_ ) );
BUF_X4 _08121_ ( .A(_01051_ ), .Z(_01052_ ) );
BUF_X4 _08122_ ( .A(_01052_ ), .Z(_01053_ ) );
BUF_X4 _08123_ ( .A(_01053_ ), .Z(_01054_ ) );
AND2_X1 _08124_ ( .A1(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A2(\u_idu.imm_auipc_lui[13] ), .ZN(_01055_ ) );
OAI21_X1 _08125_ ( .A(_00734_ ), .B1(_00651_ ), .B2(_01055_ ), .ZN(_01056_ ) );
INV_X1 _08126_ ( .A(_00644_ ), .ZN(_01057_ ) );
AOI21_X1 _08127_ ( .A(_00925_ ), .B1(_00656_ ), .B2(_01057_ ), .ZN(_01058_ ) );
NOR2_X1 _08128_ ( .A1(_01058_ ), .A2(_00694_ ), .ZN(_01059_ ) );
AOI211_X1 _08129_ ( .A(_00898_ ), .B(_01054_ ), .C1(_01056_ ), .C2(_01059_ ), .ZN(_00122_ ) );
BUF_X4 _08130_ ( .A(_00895_ ), .Z(_01060_ ) );
BUF_X2 _08131_ ( .A(_01060_ ), .Z(_01061_ ) );
BUF_X2 _08132_ ( .A(_01024_ ), .Z(_01062_ ) );
CLKBUF_X2 _08133_ ( .A(_01062_ ), .Z(_01063_ ) );
CLKBUF_X2 _08134_ ( .A(_01063_ ), .Z(_01064_ ) );
BUF_X2 _08135_ ( .A(_01049_ ), .Z(_01065_ ) );
CLKBUF_X3 _08136_ ( .A(_01065_ ), .Z(_01066_ ) );
CLKBUF_X2 _08137_ ( .A(_01066_ ), .Z(_01067_ ) );
AOI21_X1 _08138_ ( .A(_00925_ ), .B1(_00650_ ), .B2(_00661_ ), .ZN(_01068_ ) );
AND2_X1 _08139_ ( .A1(_00700_ ), .A2(_00703_ ), .ZN(_01069_ ) );
NOR2_X1 _08140_ ( .A1(_00677_ ), .A2(\u_idu.imm_auipc_lui[14] ), .ZN(_01070_ ) );
OAI211_X1 _08141_ ( .A(_00665_ ), .B(_00732_ ), .C1(_01070_ ), .C2(_00685_ ), .ZN(_01071_ ) );
OAI21_X1 _08142_ ( .A(\u_idu.imm_auipc_lui[13] ), .B1(_00647_ ), .B2(\u_idu.imm_auipc_lui[12] ), .ZN(_01072_ ) );
AOI21_X1 _08143_ ( .A(_01071_ ), .B1(_00682_ ), .B2(_01072_ ), .ZN(_01073_ ) );
OR4_X1 _08144_ ( .A1(_00694_ ), .A2(_01068_ ), .A3(_01069_ ), .A4(_01073_ ), .ZN(_01074_ ) );
AND4_X1 _08145_ ( .A1(_01061_ ), .A2(_01064_ ), .A3(_01067_ ), .A4(_01074_ ), .ZN(_00123_ ) );
BUF_X4 _08146_ ( .A(_00896_ ), .Z(_01075_ ) );
BUF_X4 _08147_ ( .A(_01075_ ), .Z(_01076_ ) );
BUF_X4 _08148_ ( .A(_01050_ ), .Z(_01077_ ) );
BUF_X2 _08149_ ( .A(_01077_ ), .Z(_01078_ ) );
AND3_X1 _08150_ ( .A1(_00700_ ), .A2(_00647_ ), .A3(_00651_ ), .ZN(_01079_ ) );
AOI21_X1 _08151_ ( .A(_01079_ ), .B1(_00727_ ), .B2(_00740_ ), .ZN(_01080_ ) );
AND3_X2 _08152_ ( .A1(_01080_ ), .A2(_00674_ ), .A3(_00747_ ), .ZN(_01081_ ) );
AND2_X1 _08153_ ( .A1(_00719_ ), .A2(_00732_ ), .ZN(_01082_ ) );
INV_X1 _08154_ ( .A(_01082_ ), .ZN(_01083_ ) );
NAND2_X1 _08155_ ( .A1(_01081_ ), .A2(_01083_ ), .ZN(_01084_ ) );
NAND3_X1 _08156_ ( .A1(_00642_ ), .A2(_00648_ ), .A3(_00657_ ), .ZN(_01085_ ) );
AND2_X1 _08157_ ( .A1(_01085_ ), .A2(_00659_ ), .ZN(_01086_ ) );
AOI21_X1 _08158_ ( .A(_00925_ ), .B1(_01086_ ), .B2(_00654_ ), .ZN(_01087_ ) );
OAI21_X1 _08159_ ( .A(\u_idu.imm_auipc_lui[14] ), .B1(_00651_ ), .B2(_00657_ ), .ZN(_01088_ ) );
OAI21_X1 _08160_ ( .A(_01088_ ), .B1(_01070_ ), .B2(_00685_ ), .ZN(_01089_ ) );
NAND2_X1 _08161_ ( .A1(_01089_ ), .A2(_00734_ ), .ZN(_01090_ ) );
NOR2_X1 _08162_ ( .A1(_00684_ ), .A2(_00687_ ), .ZN(_01091_ ) );
OAI21_X1 _08163_ ( .A(_01090_ ), .B1(_00693_ ), .B2(_01091_ ), .ZN(_01092_ ) );
NOR3_X1 _08164_ ( .A1(_01084_ ), .A2(_01087_ ), .A3(_01092_ ), .ZN(_01093_ ) );
AOI21_X1 _08165_ ( .A(_01076_ ), .B1(_01078_ ), .B2(_01093_ ), .ZN(_00124_ ) );
NOR2_X1 _08166_ ( .A1(_00742_ ), .A2(_00673_ ), .ZN(_01094_ ) );
AOI21_X1 _08167_ ( .A(_00897_ ), .B1(_00759_ ), .B2(_01094_ ), .ZN(_00231_ ) );
OAI21_X1 _08168_ ( .A(_00727_ ), .B1(_00703_ ), .B2(_00687_ ), .ZN(_01095_ ) );
OAI21_X1 _08169_ ( .A(_00671_ ), .B1(_00703_ ), .B2(_00657_ ), .ZN(_01096_ ) );
INV_X1 _08170_ ( .A(_00705_ ), .ZN(_01097_ ) );
AND3_X1 _08171_ ( .A1(_01095_ ), .A2(_01096_ ), .A3(_01097_ ), .ZN(_01098_ ) );
NAND4_X1 _08172_ ( .A1(_00700_ ), .A2(_00753_ ), .A3(_00755_ ), .A4(_00752_ ), .ZN(_01099_ ) );
NOR2_X1 _08173_ ( .A1(_01099_ ), .A2(_00715_ ), .ZN(_01100_ ) );
INV_X1 _08174_ ( .A(_01100_ ), .ZN(_01101_ ) );
OAI22_X1 _08175_ ( .A1(_00727_ ), .A2(_00700_ ), .B1(_00684_ ), .B2(_00703_ ), .ZN(_01102_ ) );
AND2_X1 _08176_ ( .A1(_01101_ ), .A2(_01102_ ), .ZN(_01103_ ) );
OAI211_X1 _08177_ ( .A(_00670_ ), .B(_00665_ ), .C1(_00703_ ), .C2(_00651_ ), .ZN(_01104_ ) );
AND2_X1 _08178_ ( .A1(_01103_ ), .A2(_01104_ ), .ZN(_01105_ ) );
AND4_X1 _08179_ ( .A1(_01078_ ), .A2(_00231_ ), .A3(_01098_ ), .A4(_01105_ ), .ZN(_00125_ ) );
OAI21_X1 _08180_ ( .A(_00692_ ), .B1(_00680_ ), .B2(_00684_ ), .ZN(_01106_ ) );
AND2_X1 _08181_ ( .A1(_00886_ ), .A2(_00713_ ), .ZN(_01107_ ) );
AND4_X1 _08182_ ( .A1(_00751_ ), .A2(_00638_ ), .A3(_00641_ ), .A4(_00711_ ), .ZN(_01108_ ) );
NAND3_X1 _08183_ ( .A1(_01108_ ), .A2(_00893_ ), .A3(_00753_ ), .ZN(_01109_ ) );
NAND2_X1 _08184_ ( .A1(_00756_ ), .A2(_01109_ ), .ZN(_01110_ ) );
OAI21_X1 _08185_ ( .A(_00686_ ), .B1(_01107_ ), .B2(_01110_ ), .ZN(_01111_ ) );
AOI21_X1 _08186_ ( .A(_00701_ ), .B1(_01111_ ), .B2(_00704_ ), .ZN(_01112_ ) );
NOR2_X1 _08187_ ( .A1(_01112_ ), .A2(_00698_ ), .ZN(_01113_ ) );
AOI211_X1 _08188_ ( .A(_00766_ ), .B(_00874_ ), .C1(_01106_ ), .C2(_01113_ ), .ZN(_00229_ ) );
AND3_X1 _08189_ ( .A1(_01064_ ), .A2(_01067_ ), .A3(_00229_ ), .ZN(_00126_ ) );
OR2_X1 _08190_ ( .A1(_00693_ ), .A2(_01088_ ), .ZN(_01114_ ) );
NOR2_X1 _08191_ ( .A1(_00862_ ), .A2(\u_idu.imm_auipc_lui[31] ), .ZN(_01115_ ) );
NAND2_X1 _08192_ ( .A1(_00652_ ), .A2(_01115_ ), .ZN(_01116_ ) );
NAND3_X1 _08193_ ( .A1(_00646_ ), .A2(_00640_ ), .A3(_00643_ ), .ZN(_01117_ ) );
NAND2_X1 _08194_ ( .A1(_01116_ ), .A2(_01117_ ), .ZN(_01118_ ) );
NAND2_X1 _08195_ ( .A1(_01118_ ), .A2(_00668_ ), .ZN(_01119_ ) );
OAI21_X1 _08196_ ( .A(_00671_ ), .B1(_00684_ ), .B2(_00687_ ), .ZN(_01120_ ) );
INV_X1 _08197_ ( .A(\u_exu.opt_$_NOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B ), .ZN(_01121_ ) );
AND4_X1 _08198_ ( .A1(\u_idu.imm_auipc_lui[12] ), .A2(_00677_ ), .A3(_01121_ ), .A4(\u_idu.imm_auipc_lui[14] ), .ZN(_01122_ ) );
OAI21_X1 _08199_ ( .A(_00734_ ), .B1(_00703_ ), .B2(_01122_ ), .ZN(_01123_ ) );
AND3_X1 _08200_ ( .A1(_01119_ ), .A2(_01120_ ), .A3(_01123_ ), .ZN(_01124_ ) );
AOI211_X1 _08201_ ( .A(_00766_ ), .B(_00874_ ), .C1(_01114_ ), .C2(_01124_ ), .ZN(_00230_ ) );
AND3_X1 _08202_ ( .A1(_01064_ ), .A2(_01067_ ), .A3(_00230_ ), .ZN(_00127_ ) );
OAI21_X1 _08203_ ( .A(_00734_ ), .B1(_01070_ ), .B2(_00681_ ), .ZN(_01125_ ) );
NAND2_X1 _08204_ ( .A1(_00658_ ), .A2(_01115_ ), .ZN(_01126_ ) );
AOI21_X1 _08205_ ( .A(_00925_ ), .B1(_00650_ ), .B2(_01126_ ), .ZN(_01127_ ) );
NOR3_X1 _08206_ ( .A1(_01127_ ), .A2(_00694_ ), .A3(_01069_ ), .ZN(_01128_ ) );
AOI211_X1 _08207_ ( .A(_00898_ ), .B(_01054_ ), .C1(_01125_ ), .C2(_01128_ ), .ZN(_00128_ ) );
INV_X1 _08208_ ( .A(fanout_net_11 ), .ZN(_01129_ ) );
INV_X32 _08209_ ( .A(icah_valid ), .ZN(_01130_ ) );
NOR2_X4 _08210_ ( .A1(_01130_ ), .A2(\u_arbiter.working ), .ZN(_01131_ ) );
BUF_X4 _08211_ ( .A(_01131_ ), .Z(_01132_ ) );
NAND2_X1 _08212_ ( .A1(_01132_ ), .A2(io_master_rready_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A ), .ZN(_01133_ ) );
BUF_X4 _08213_ ( .A(_01130_ ), .Z(_01134_ ) );
OAI21_X1 _08214_ ( .A(io_master_rready_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_MUX__Y_B ), .B1(_01134_ ), .B2(\u_arbiter.working ), .ZN(_01135_ ) );
AND2_X1 _08215_ ( .A1(_01133_ ), .A2(_01135_ ), .ZN(_01136_ ) );
BUF_X4 _08216_ ( .A(_01132_ ), .Z(_01137_ ) );
NOR2_X1 _08217_ ( .A1(_01137_ ), .A2(\u_arbiter.raddr[11] ), .ZN(_01138_ ) );
NOR3_X1 _08218_ ( .A1(_01134_ ), .A2(\u_arbiter.working ), .A3(\ca_addr[11] ), .ZN(_01139_ ) );
NOR2_X1 _08219_ ( .A1(_01138_ ), .A2(_01139_ ), .ZN(\io_master_araddr[11] ) );
OR2_X1 _08220_ ( .A1(_01136_ ), .A2(\io_master_araddr[11] ), .ZN(_01140_ ) );
BUF_X4 _08221_ ( .A(_01132_ ), .Z(_01141_ ) );
NAND2_X1 _08222_ ( .A1(_01141_ ), .A2(\ca_addr[15] ), .ZN(_01142_ ) );
BUF_X4 _08223_ ( .A(_01134_ ), .Z(_01143_ ) );
OAI21_X1 _08224_ ( .A(\u_arbiter.raddr[15] ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_01144_ ) );
NAND2_X1 _08225_ ( .A1(_01142_ ), .A2(_01144_ ), .ZN(\io_master_araddr[15] ) );
NAND2_X1 _08226_ ( .A1(_01141_ ), .A2(\ca_addr[12] ), .ZN(_01145_ ) );
OAI21_X1 _08227_ ( .A(\u_arbiter.raddr[12] ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_01146_ ) );
NAND2_X1 _08228_ ( .A1(_01145_ ), .A2(_01146_ ), .ZN(\io_master_araddr[12] ) );
NOR3_X1 _08229_ ( .A1(_01140_ ), .A2(\io_master_araddr[15] ), .A3(\io_master_araddr[12] ), .ZN(_01147_ ) );
MUX2_X1 _08230_ ( .A(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_B ), .B(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_A ), .S(_01131_ ), .Z(_01148_ ) );
INV_X1 _08231_ ( .A(_01148_ ), .ZN(\io_master_araddr[10] ) );
MUX2_X1 _08232_ ( .A(\u_arbiter.raddr[13] ), .B(\ca_addr[13] ), .S(_01132_ ), .Z(\io_master_araddr[13] ) );
OR2_X1 _08233_ ( .A1(\io_master_araddr[10] ), .A2(\io_master_araddr[13] ), .ZN(_01149_ ) );
MUX2_X1 _08234_ ( .A(\u_arbiter.raddr[14] ), .B(\ca_addr[14] ), .S(_01137_ ), .Z(\io_master_araddr[14] ) );
MUX2_X1 _08235_ ( .A(\u_arbiter.raddr[9] ), .B(\ca_addr[9] ), .S(_01137_ ), .Z(\io_master_araddr[9] ) );
NOR3_X2 _08236_ ( .A1(_01149_ ), .A2(\io_master_araddr[14] ), .A3(\io_master_araddr[9] ), .ZN(_01150_ ) );
NAND2_X1 _08237_ ( .A1(_01141_ ), .A2(\ca_addr[17] ), .ZN(_01151_ ) );
NAND2_X1 _08238_ ( .A1(_01137_ ), .A2(\ca_addr[22] ), .ZN(_01152_ ) );
OAI21_X1 _08239_ ( .A(\u_arbiter.raddr[17] ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_01153_ ) );
OAI21_X1 _08240_ ( .A(\u_arbiter.raddr[22] ), .B1(_01134_ ), .B2(\u_arbiter.working ), .ZN(_01154_ ) );
NAND4_X1 _08241_ ( .A1(_01151_ ), .A2(_01152_ ), .A3(_01153_ ), .A4(_01154_ ), .ZN(_01155_ ) );
NAND2_X1 _08242_ ( .A1(_01137_ ), .A2(\ca_addr[18] ), .ZN(_01156_ ) );
NAND2_X1 _08243_ ( .A1(_01137_ ), .A2(\ca_addr[21] ), .ZN(_01157_ ) );
OAI21_X1 _08244_ ( .A(\u_arbiter.raddr[18] ), .B1(_01134_ ), .B2(\u_arbiter.working ), .ZN(_01158_ ) );
OAI21_X1 _08245_ ( .A(\u_arbiter.raddr[21] ), .B1(_01134_ ), .B2(\u_arbiter.working ), .ZN(_01159_ ) );
NAND4_X1 _08246_ ( .A1(_01156_ ), .A2(_01157_ ), .A3(_01158_ ), .A4(_01159_ ), .ZN(_01160_ ) );
NOR2_X1 _08247_ ( .A1(_01155_ ), .A2(_01160_ ), .ZN(_01161_ ) );
MUX2_X1 _08248_ ( .A(\u_arbiter.raddr[26] ), .B(\ca_addr[26] ), .S(_01132_ ), .Z(\io_master_araddr[26] ) );
NAND2_X1 _08249_ ( .A1(_01137_ ), .A2(\ca_addr[27] ), .ZN(_01162_ ) );
OAI21_X1 _08250_ ( .A(\u_arbiter.raddr[27] ), .B1(_01134_ ), .B2(\u_arbiter.working ), .ZN(_01163_ ) );
NAND2_X1 _08251_ ( .A1(_01162_ ), .A2(_01163_ ), .ZN(\io_master_araddr[27] ) );
NOR2_X1 _08252_ ( .A1(\io_master_araddr[26] ), .A2(\io_master_araddr[27] ), .ZN(_01164_ ) );
OR3_X1 _08253_ ( .A1(_01134_ ), .A2(\u_arbiter.working ), .A3(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_A ), .ZN(_01165_ ) );
OAI21_X1 _08254_ ( .A(_01165_ ), .B1(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_B ), .B2(_01137_ ), .ZN(\io_master_araddr[25] ) );
NAND2_X1 _08255_ ( .A1(_01137_ ), .A2(\ca_addr[24] ), .ZN(_01166_ ) );
OAI21_X1 _08256_ ( .A(\u_arbiter.raddr[24] ), .B1(_01134_ ), .B2(\u_arbiter.working ), .ZN(_01167_ ) );
NAND2_X1 _08257_ ( .A1(_01166_ ), .A2(_01167_ ), .ZN(\io_master_araddr[24] ) );
NOR2_X1 _08258_ ( .A1(\io_master_araddr[25] ), .A2(\io_master_araddr[24] ), .ZN(_01168_ ) );
AND2_X1 _08259_ ( .A1(_01164_ ), .A2(_01168_ ), .ZN(_01169_ ) );
AND3_X1 _08260_ ( .A1(_01150_ ), .A2(_01161_ ), .A3(_01169_ ), .ZN(_01170_ ) );
MUX2_X1 _08261_ ( .A(\u_arbiter.raddr[19] ), .B(\ca_addr[19] ), .S(_01141_ ), .Z(\io_master_araddr[19] ) );
MUX2_X1 _08262_ ( .A(\u_arbiter.raddr[23] ), .B(\ca_addr[23] ), .S(_01137_ ), .Z(\io_master_araddr[23] ) );
NOR2_X1 _08263_ ( .A1(\io_master_araddr[19] ), .A2(\io_master_araddr[23] ), .ZN(_01171_ ) );
NOR2_X1 _08264_ ( .A1(_01141_ ), .A2(\u_arbiter.raddr[20] ), .ZN(_01172_ ) );
NOR3_X1 _08265_ ( .A1(_01143_ ), .A2(\u_arbiter.working ), .A3(\ca_addr[20] ), .ZN(_01173_ ) );
NOR2_X1 _08266_ ( .A1(_01172_ ), .A2(_01173_ ), .ZN(\io_master_araddr[20] ) );
NAND2_X1 _08267_ ( .A1(_01141_ ), .A2(\ca_addr[16] ), .ZN(_01174_ ) );
OAI21_X1 _08268_ ( .A(\u_arbiter.raddr[16] ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_01175_ ) );
NAND2_X1 _08269_ ( .A1(_01174_ ), .A2(_01175_ ), .ZN(\io_master_araddr[16] ) );
NOR2_X1 _08270_ ( .A1(\io_master_araddr[20] ), .A2(\io_master_araddr[16] ), .ZN(_01176_ ) );
AND4_X2 _08271_ ( .A1(_01147_ ), .A2(_01170_ ), .A3(_01171_ ), .A4(_01176_ ), .ZN(_01177_ ) );
NAND2_X1 _08272_ ( .A1(_01131_ ), .A2(\ca_addr[7] ), .ZN(_01178_ ) );
OAI21_X1 _08273_ ( .A(\u_arbiter.raddr[7] ), .B1(_01134_ ), .B2(\u_arbiter.working ), .ZN(_01179_ ) );
NAND2_X1 _08274_ ( .A1(_01178_ ), .A2(_01179_ ), .ZN(\io_master_araddr[7] ) );
INV_X1 _08275_ ( .A(\io_master_araddr[7] ), .ZN(_01180_ ) );
MUX2_X1 _08276_ ( .A(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_B ), .B(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_A ), .S(_01132_ ), .Z(_01181_ ) );
INV_X1 _08277_ ( .A(_01181_ ), .ZN(\io_master_araddr[4] ) );
MUX2_X1 _08278_ ( .A(\u_arbiter.raddr[5] ), .B(\ca_addr[5] ), .S(_01132_ ), .Z(\io_master_araddr[5] ) );
NOR2_X1 _08279_ ( .A1(\io_master_araddr[4] ), .A2(\io_master_araddr[5] ), .ZN(_01182_ ) );
OR3_X4 _08280_ ( .A1(_01130_ ), .A2(\u_arbiter.working ), .A3(io_master_araddr_$_NOT__Y_A_$_MUX__Y_A ), .ZN(_01183_ ) );
OAI21_X1 _08281_ ( .A(_01183_ ), .B1(io_master_araddr_$_NOT__Y_A_$_MUX__Y_B ), .B2(_01132_ ), .ZN(\io_master_araddr[6] ) );
AND2_X1 _08282_ ( .A1(_01180_ ), .A2(\io_master_araddr[6] ), .ZN(_01184_ ) );
INV_X1 _08283_ ( .A(_01184_ ), .ZN(_01185_ ) );
OAI211_X1 _08284_ ( .A(_01177_ ), .B(_01180_ ), .C1(_01182_ ), .C2(_01185_ ), .ZN(_01186_ ) );
NOR2_X1 _08285_ ( .A1(_01141_ ), .A2(\u_arbiter.raddr[31] ), .ZN(_01187_ ) );
NOR3_X1 _08286_ ( .A1(_01143_ ), .A2(\u_arbiter.working ), .A3(\ca_addr[31] ), .ZN(_01188_ ) );
NOR2_X1 _08287_ ( .A1(_01187_ ), .A2(_01188_ ), .ZN(\io_master_araddr[31] ) );
NAND2_X1 _08288_ ( .A1(_01141_ ), .A2(\ca_addr[29] ), .ZN(_01189_ ) );
OAI21_X1 _08289_ ( .A(\u_arbiter.raddr[29] ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_01190_ ) );
NAND2_X1 _08290_ ( .A1(_01189_ ), .A2(_01190_ ), .ZN(\io_master_araddr[29] ) );
AND2_X1 _08291_ ( .A1(\io_master_araddr[31] ), .A2(\io_master_araddr[29] ), .ZN(_01191_ ) );
NAND2_X2 _08292_ ( .A1(_01186_ ), .A2(_01191_ ), .ZN(_01192_ ) );
NAND2_X1 _08293_ ( .A1(_01141_ ), .A2(\ca_addr[30] ), .ZN(_01193_ ) );
OAI21_X1 _08294_ ( .A(\u_arbiter.raddr[30] ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_01194_ ) );
NAND2_X1 _08295_ ( .A1(_01193_ ), .A2(_01194_ ), .ZN(\io_master_araddr[30] ) );
BUF_X2 _08296_ ( .A(_01141_ ), .Z(_01195_ ) );
NAND2_X1 _08297_ ( .A1(_01195_ ), .A2(\ca_addr[28] ), .ZN(_01196_ ) );
OAI21_X1 _08298_ ( .A(\u_arbiter.raddr[28] ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_01197_ ) );
NAND2_X1 _08299_ ( .A1(_01196_ ), .A2(_01197_ ), .ZN(\io_master_araddr[28] ) );
INV_X1 _08300_ ( .A(_01132_ ), .ZN(_01198_ ) );
AND2_X1 _08301_ ( .A1(_01198_ ), .A2(\u_arbiter.raddr[3] ), .ZN(_01199_ ) );
NOR3_X1 _08302_ ( .A1(\io_master_araddr[4] ), .A2(\io_master_araddr[5] ), .A3(_01199_ ), .ZN(_01200_ ) );
MUX2_X1 _08303_ ( .A(\u_arbiter.raddr[8] ), .B(\ca_addr[8] ), .S(_01132_ ), .Z(\io_master_araddr[8] ) );
OR3_X4 _08304_ ( .A1(_01200_ ), .A2(_01185_ ), .A3(\io_master_araddr[8] ), .ZN(_01201_ ) );
NAND4_X1 _08305_ ( .A1(_01201_ ), .A2(_01180_ ), .A3(_01171_ ), .A4(_01176_ ), .ZN(_01202_ ) );
NAND4_X1 _08306_ ( .A1(_01150_ ), .A2(_01147_ ), .A3(_01161_ ), .A4(_01169_ ), .ZN(_01203_ ) );
OAI221_X1 _08307_ ( .A(\io_master_araddr[31] ), .B1(\io_master_araddr[29] ), .B2(\io_master_araddr[30] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_01204_ ) );
BUF_X4 _08308_ ( .A(_01198_ ), .Z(_01205_ ) );
INV_X1 _08309_ ( .A(\u_arbiter.raddr[0] ), .ZN(_01206_ ) );
INV_X1 _08310_ ( .A(\u_arbiter.raddr[1] ), .ZN(_01207_ ) );
NAND4_X4 _08311_ ( .A1(_01205_ ), .A2(\u_arbiter.raddr[3] ), .A3(_01206_ ), .A4(_01207_ ), .ZN(_01208_ ) );
NOR2_X2 _08312_ ( .A1(_01208_ ), .A2(\u_arbiter.raddr[2] ), .ZN(_01209_ ) );
NAND4_X1 _08313_ ( .A1(_01182_ ), .A2(_01191_ ), .A3(_01184_ ), .A4(_01209_ ), .ZN(_01210_ ) );
AOI211_X2 _08314_ ( .A(\io_master_araddr[30] ), .B(\io_master_araddr[28] ), .C1(_01204_ ), .C2(_01210_ ), .ZN(_01211_ ) );
AND2_X4 _08315_ ( .A1(_01192_ ), .A2(_01211_ ), .ZN(_01212_ ) );
AND2_X4 _08316_ ( .A1(_01212_ ), .A2(\u_lsu.rvalid_clint ), .ZN(_01213_ ) );
INV_X1 _08317_ ( .A(_01212_ ), .ZN(_01214_ ) );
AOI21_X4 _08318_ ( .A(_01213_ ), .B1(io_master_rvalid ), .B2(_01214_ ), .ZN(_01215_ ) );
INV_X1 _08319_ ( .A(\u_lsu.reading ), .ZN(_01216_ ) );
MUX2_X1 _08320_ ( .A(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_A ), .B(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ), .S(_01195_ ), .Z(_01217_ ) );
OR4_X2 _08321_ ( .A1(_01129_ ), .A2(_01215_ ), .A3(_01216_ ), .A4(_01217_ ), .ZN(_01218_ ) );
AOI211_X1 _08322_ ( .A(ea_err ), .B(_00763_ ), .C1(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ), .C2(_00629_ ), .ZN(_01219_ ) );
NAND2_X1 _08323_ ( .A1(_01219_ ), .A2(\u_exu.eopt[0] ), .ZN(_01220_ ) );
AND2_X4 _08324_ ( .A1(_01218_ ), .A2(_01220_ ), .ZN(_01221_ ) );
BUF_X4 _08325_ ( .A(_01221_ ), .Z(_01222_ ) );
INV_X4 _08326_ ( .A(_01222_ ), .ZN(_01223_ ) );
NAND2_X1 _08327_ ( .A1(_01129_ ), .A2(\ea_ard[0] ), .ZN(_01224_ ) );
NAND2_X1 _08328_ ( .A1(fanout_net_11 ), .A2(\u_arbiter.wbaddr[0] ), .ZN(_01225_ ) );
NAND2_X1 _08329_ ( .A1(_01224_ ), .A2(_01225_ ), .ZN(_01226_ ) );
XNOR2_X1 _08330_ ( .A(_00904_ ), .B(_01226_ ), .ZN(_01227_ ) );
NAND2_X1 _08331_ ( .A1(_01129_ ), .A2(\ea_ard[3] ), .ZN(_01228_ ) );
NAND2_X1 _08332_ ( .A1(\u_arbiter.wbaddr[3] ), .A2(fanout_net_11 ), .ZN(_01229_ ) );
NAND2_X1 _08333_ ( .A1(_01228_ ), .A2(_01229_ ), .ZN(_01230_ ) );
INV_X2 _08334_ ( .A(_01230_ ), .ZN(_01231_ ) );
XNOR2_X1 _08335_ ( .A(_00912_ ), .B(_01231_ ), .ZN(_01232_ ) );
NAND2_X1 _08336_ ( .A1(_01129_ ), .A2(\ea_ard[1] ), .ZN(_01233_ ) );
NAND2_X1 _08337_ ( .A1(fanout_net_11 ), .A2(\u_arbiter.wbaddr[1] ), .ZN(_01234_ ) );
NAND2_X1 _08338_ ( .A1(_01233_ ), .A2(_01234_ ), .ZN(_01235_ ) );
XNOR2_X1 _08339_ ( .A(_00907_ ), .B(_01235_ ), .ZN(_01236_ ) );
NAND2_X1 _08340_ ( .A1(_01129_ ), .A2(\ea_ard[2] ), .ZN(_01237_ ) );
NAND2_X1 _08341_ ( .A1(fanout_net_11 ), .A2(\u_arbiter.wbaddr[2] ), .ZN(_01238_ ) );
NAND2_X2 _08342_ ( .A1(_01237_ ), .A2(_01238_ ), .ZN(_01239_ ) );
INV_X1 _08343_ ( .A(_01239_ ), .ZN(_01240_ ) );
NAND3_X1 _08344_ ( .A1(_00902_ ), .A2(_00913_ ), .A3(_01240_ ), .ZN(_01241_ ) );
NAND4_X1 _08345_ ( .A1(_01227_ ), .A2(_01232_ ), .A3(_01236_ ), .A4(_01241_ ), .ZN(_01242_ ) );
AOI21_X1 _08346_ ( .A(_01242_ ), .B1(_00975_ ), .B2(_01239_ ), .ZN(_01243_ ) );
AND2_X2 _08347_ ( .A1(_01223_ ), .A2(_01243_ ), .ZN(_01244_ ) );
INV_X1 _08348_ ( .A(_01244_ ), .ZN(_01245_ ) );
BUF_X4 _08349_ ( .A(_01245_ ), .Z(_01246_ ) );
NOR2_X1 _08350_ ( .A1(_01209_ ), .A2(\u_lsu.u_clint.mtime[47] ), .ZN(_01247_ ) );
INV_X1 _08351_ ( .A(_01213_ ), .ZN(_01248_ ) );
INV_X1 _08352_ ( .A(\u_lsu.u_clint.mtime[15] ), .ZN(_01249_ ) );
AOI211_X2 _08353_ ( .A(_01247_ ), .B(_01248_ ), .C1(_01249_ ), .C2(_01209_ ), .ZN(_01250_ ) );
AOI21_X1 _08354_ ( .A(_01250_ ), .B1(_01214_ ), .B2(\io_master_rdata[15] ), .ZN(_01251_ ) );
NOR2_X1 _08355_ ( .A1(_01195_ ), .A2(_01207_ ), .ZN(\io_master_araddr[1] ) );
NOR2_X1 _08356_ ( .A1(_01195_ ), .A2(_01206_ ), .ZN(\io_master_araddr[0] ) );
NOR2_X1 _08357_ ( .A1(\io_master_araddr[1] ), .A2(\io_master_araddr[0] ), .ZN(_01252_ ) );
INV_X1 _08358_ ( .A(_01252_ ), .ZN(_01253_ ) );
OR2_X1 _08359_ ( .A1(_01251_ ), .A2(_01253_ ), .ZN(_01254_ ) );
AND2_X2 _08360_ ( .A1(\io_master_araddr[1] ), .A2(_01206_ ), .ZN(_01255_ ) );
INV_X1 _08361_ ( .A(_01255_ ), .ZN(_01256_ ) );
INV_X1 _08362_ ( .A(\u_arbiter.raddr[2] ), .ZN(_01257_ ) );
BUF_X4 _08363_ ( .A(_01257_ ), .Z(_01258_ ) );
BUF_X2 _08364_ ( .A(_01199_ ), .Z(\io_master_araddr[3] ) );
INV_X1 _08365_ ( .A(\u_lsu.u_clint.mtime[31] ), .ZN(_01259_ ) );
NAND4_X1 _08366_ ( .A1(_01252_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_01259_ ), .ZN(_01260_ ) );
OAI211_X1 _08367_ ( .A(_01213_ ), .B(_01260_ ), .C1(\u_lsu.u_clint.mtime[63] ), .C2(_01209_ ), .ZN(_01261_ ) );
NAND2_X1 _08368_ ( .A1(_01214_ ), .A2(\io_master_rdata[31] ), .ZN(_01262_ ) );
AOI21_X1 _08369_ ( .A(_01256_ ), .B1(_01261_ ), .B2(_01262_ ), .ZN(_01263_ ) );
INV_X1 _08370_ ( .A(\u_lsu.u_clint.mtime[23] ), .ZN(_01264_ ) );
NAND4_X1 _08371_ ( .A1(_01252_ ), .A2(_01257_ ), .A3(_01199_ ), .A4(_01264_ ), .ZN(_01265_ ) );
OAI211_X1 _08372_ ( .A(_01213_ ), .B(_01265_ ), .C1(\u_lsu.u_clint.mtime[55] ), .C2(_01209_ ), .ZN(_01266_ ) );
NAND2_X1 _08373_ ( .A1(_01214_ ), .A2(\io_master_rdata[23] ), .ZN(_01267_ ) );
AND2_X1 _08374_ ( .A1(_01266_ ), .A2(_01267_ ), .ZN(_01268_ ) );
INV_X1 _08375_ ( .A(_01268_ ), .ZN(_01269_ ) );
AND2_X2 _08376_ ( .A1(\io_master_araddr[0] ), .A2(_01207_ ), .ZN(_01270_ ) );
AOI21_X1 _08377_ ( .A(_01263_ ), .B1(_01269_ ), .B2(_01270_ ), .ZN(_01271_ ) );
AND2_X1 _08378_ ( .A1(_01254_ ), .A2(_01271_ ), .ZN(_01272_ ) );
NOR2_X1 _08379_ ( .A1(_01195_ ), .A2(\u_arbiter.rmask[0] ), .ZN(_01273_ ) );
NAND3_X1 _08380_ ( .A1(_01273_ ), .A2(\u_arbiter.rmask[1] ), .A3(\u_arbiter.rsign ), .ZN(_01274_ ) );
NOR2_X4 _08381_ ( .A1(_01272_ ), .A2(_01274_ ), .ZN(_01275_ ) );
BUF_X2 _08382_ ( .A(_01252_ ), .Z(_01276_ ) );
NOR2_X1 _08383_ ( .A1(_01195_ ), .A2(\u_arbiter.rmask[1] ), .ZN(_01277_ ) );
NOR2_X1 _08384_ ( .A1(_01277_ ), .A2(_01273_ ), .ZN(_01278_ ) );
NAND2_X1 _08385_ ( .A1(_01276_ ), .A2(_01278_ ), .ZN(_01279_ ) );
AOI21_X1 _08386_ ( .A(_01279_ ), .B1(_01261_ ), .B2(_01262_ ), .ZN(_01280_ ) );
AND2_X1 _08387_ ( .A1(\io_master_araddr[1] ), .A2(\u_arbiter.raddr[0] ), .ZN(_01281_ ) );
INV_X1 _08388_ ( .A(_01281_ ), .ZN(_01282_ ) );
AOI21_X1 _08389_ ( .A(_01282_ ), .B1(_01261_ ), .B2(_01262_ ), .ZN(_01283_ ) );
AOI21_X1 _08390_ ( .A(_01283_ ), .B1(_01269_ ), .B2(_01255_ ), .ZN(_01284_ ) );
INV_X1 _08391_ ( .A(_01270_ ), .ZN(_01285_ ) );
OAI21_X1 _08392_ ( .A(_01284_ ), .B1(_01251_ ), .B2(_01285_ ), .ZN(_01286_ ) );
NAND2_X1 _08393_ ( .A1(_01214_ ), .A2(\io_master_rdata[7] ), .ZN(_01287_ ) );
MUX2_X1 _08394_ ( .A(\u_lsu.u_clint.mtime[39] ), .B(\u_lsu.u_clint.mtime[7] ), .S(_01209_ ), .Z(_01288_ ) );
NAND4_X1 _08395_ ( .A1(_01192_ ), .A2(_01211_ ), .A3(\u_lsu.rvalid_clint ), .A4(_01288_ ), .ZN(_01289_ ) );
AOI21_X1 _08396_ ( .A(_01253_ ), .B1(_01287_ ), .B2(_01289_ ), .ZN(_01290_ ) );
NOR2_X2 _08397_ ( .A1(_01286_ ), .A2(_01290_ ), .ZN(_01291_ ) );
INV_X1 _08398_ ( .A(\u_arbiter.rmask[1] ), .ZN(_01292_ ) );
NAND4_X1 _08399_ ( .A1(_01205_ ), .A2(_01292_ ), .A3(\u_arbiter.rmask[0] ), .A4(\u_arbiter.rsign ), .ZN(_01293_ ) );
NOR2_X2 _08400_ ( .A1(_01291_ ), .A2(_01293_ ), .ZN(_01294_ ) );
BUF_X4 _08401_ ( .A(_01294_ ), .Z(_01295_ ) );
NOR3_X1 _08402_ ( .A1(_01275_ ), .A2(_01280_ ), .A3(_01295_ ), .ZN(_01296_ ) );
NAND2_X1 _08403_ ( .A1(_01296_ ), .A2(fanout_net_11 ), .ZN(_01297_ ) );
AND2_X2 _08404_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .ZN(_01298_ ) );
BUF_X4 _08405_ ( .A(_01298_ ), .Z(_01299_ ) );
MUX2_X1 _08406_ ( .A(\ea_addr[31] ), .B(\u_exu.ecsr[31] ), .S(_01299_ ), .Z(_01300_ ) );
OR2_X1 _08407_ ( .A1(_01300_ ), .A2(fanout_net_11 ), .ZN(_01301_ ) );
AOI21_X1 _08408_ ( .A(_01246_ ), .B1(_01297_ ), .B2(_01301_ ), .ZN(_01302_ ) );
BUF_X4 _08409_ ( .A(_00736_ ), .Z(_01303_ ) );
BUF_X4 _08410_ ( .A(_01244_ ), .Z(_01304_ ) );
BUF_X4 _08411_ ( .A(_00950_ ), .Z(_01305_ ) );
BUF_X4 _08412_ ( .A(_00909_ ), .Z(_01306_ ) );
AOI22_X1 _08413_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01307_ ) );
BUF_X4 _08414_ ( .A(_01005_ ), .Z(_01308_ ) );
NOR2_X2 _08415_ ( .A1(_00904_ ), .A2(_00907_ ), .ZN(_01309_ ) );
BUF_X4 _08416_ ( .A(_01309_ ), .Z(_01310_ ) );
AOI22_X1 _08417_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01311_ ) );
BUF_X4 _08418_ ( .A(_00975_ ), .Z(_01312_ ) );
NAND3_X1 _08419_ ( .A1(_01307_ ), .A2(_01311_ ), .A3(_01312_ ), .ZN(_01313_ ) );
BUF_X4 _08420_ ( .A(_01309_ ), .Z(_01314_ ) );
AOI22_X1 _08421_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01315_ ) );
BUF_X4 _08422_ ( .A(_00950_ ), .Z(_01316_ ) );
AOI22_X1 _08423_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01317_ ) );
BUF_X2 _08424_ ( .A(_00915_ ), .Z(_01318_ ) );
NAND3_X1 _08425_ ( .A1(_01315_ ), .A2(_01317_ ), .A3(_01318_ ), .ZN(_01319_ ) );
CLKBUF_X2 _08426_ ( .A(_00951_ ), .Z(_01320_ ) );
AND3_X1 _08427_ ( .A1(_01313_ ), .A2(_01319_ ), .A3(_01320_ ), .ZN(_01321_ ) );
BUF_X4 _08428_ ( .A(_00902_ ), .Z(_01322_ ) );
BUF_X4 _08429_ ( .A(_00907_ ), .Z(_01323_ ) );
OAI211_X1 _08430_ ( .A(fanout_net_21 ), .B(_01322_ ), .C1(_01323_ ), .C2(\u_reg.rf[1][31] ), .ZN(_01324_ ) );
BUF_X2 _08431_ ( .A(_00908_ ), .Z(_01325_ ) );
OAI21_X1 _08432_ ( .A(_01324_ ), .B1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01325_ ), .ZN(_01326_ ) );
BUF_X4 _08433_ ( .A(_00975_ ), .Z(_01327_ ) );
BUF_X4 _08434_ ( .A(_01323_ ), .Z(_01328_ ) );
NAND4_X1 _08435_ ( .A1(_01328_ ), .A2(fanout_net_21 ), .A3(_01322_ ), .A4(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01329_ ) );
NAND3_X1 _08436_ ( .A1(_01326_ ), .A2(_01327_ ), .A3(_01329_ ), .ZN(_01330_ ) );
AND2_X1 _08437_ ( .A1(_01330_ ), .A2(_01046_ ), .ZN(_01331_ ) );
BUF_X4 _08438_ ( .A(_00909_ ), .Z(_01332_ ) );
BUF_X4 _08439_ ( .A(_01332_ ), .Z(_01333_ ) );
BUF_X4 _08440_ ( .A(_01310_ ), .Z(_01334_ ) );
AOI22_X1 _08441_ ( .A1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01333_ ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01335_ ) );
BUF_X4 _08442_ ( .A(_00915_ ), .Z(_01336_ ) );
BUF_X4 _08443_ ( .A(_00904_ ), .Z(_01337_ ) );
BUF_X4 _08444_ ( .A(_01337_ ), .Z(_01338_ ) );
BUF_X4 _08445_ ( .A(_01323_ ), .Z(_01339_ ) );
NAND3_X1 _08446_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01339_ ), .ZN(_01340_ ) );
BUF_X4 _08447_ ( .A(_00908_ ), .Z(_01341_ ) );
BUF_X4 _08448_ ( .A(_01341_ ), .Z(_01342_ ) );
NAND3_X1 _08449_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01342_ ), .ZN(_01343_ ) );
NAND4_X1 _08450_ ( .A1(_01335_ ), .A2(_01336_ ), .A3(_01340_ ), .A4(_01343_ ), .ZN(_01344_ ) );
AOI21_X1 _08451_ ( .A(_01321_ ), .B1(_01331_ ), .B2(_01344_ ), .ZN(_01345_ ) );
OAI21_X1 _08452_ ( .A(_01303_ ), .B1(_01304_ ), .B2(_01345_ ), .ZN(_01346_ ) );
OR3_X1 _08453_ ( .A1(_01302_ ), .A2(_00723_ ), .A3(_01346_ ), .ZN(_01347_ ) );
AND2_X1 _08454_ ( .A1(_00700_ ), .A2(_00687_ ), .ZN(_01348_ ) );
AND4_X1 _08455_ ( .A1(_00894_ ), .A2(_00709_ ), .A3(fanout_net_23 ), .A4(_00751_ ), .ZN(_01349_ ) );
AND3_X1 _08456_ ( .A1(_01349_ ), .A2(_00708_ ), .A3(_00755_ ), .ZN(_01350_ ) );
AND2_X1 _08457_ ( .A1(_01348_ ), .A2(_01350_ ), .ZN(_01351_ ) );
INV_X1 _08458_ ( .A(_01351_ ), .ZN(_01352_ ) );
BUF_X4 _08459_ ( .A(_01352_ ), .Z(_01353_ ) );
INV_X1 _08460_ ( .A(\u_exu.acsrd[11] ), .ZN(_01354_ ) );
NOR2_X1 _08461_ ( .A1(_01354_ ), .A2(ea_err ), .ZN(_01355_ ) );
NOR3_X1 _08462_ ( .A1(_00634_ ), .A2(_00653_ ), .A3(_01355_ ), .ZN(_01356_ ) );
AND2_X1 _08463_ ( .A1(_00785_ ), .A2(\u_exu.acsrd[5] ), .ZN(_01357_ ) );
INV_X1 _08464_ ( .A(_01357_ ), .ZN(_01358_ ) );
AND2_X1 _08465_ ( .A1(_00784_ ), .A2(\u_exu.acsrd[4] ), .ZN(_01359_ ) );
INV_X1 _08466_ ( .A(_01359_ ), .ZN(_01360_ ) );
AOI22_X1 _08467_ ( .A1(\u_idu.imm_auipc_lui[25] ), .A2(_01358_ ), .B1(_01360_ ), .B2(\u_idu.imm_auipc_lui[24] ), .ZN(_01361_ ) );
AND2_X1 _08468_ ( .A1(_00785_ ), .A2(\u_exu.acsrd[7] ), .ZN(_01362_ ) );
NOR2_X1 _08469_ ( .A1(ea_err ), .A2(\u_exu.acsrd[9] ), .ZN(_01363_ ) );
OAI221_X1 _08470_ ( .A(_01361_ ), .B1(_00707_ ), .B2(_01362_ ), .C1(\u_idu.imm_auipc_lui[29] ), .C2(_01363_ ), .ZN(_01364_ ) );
AOI21_X1 _08471_ ( .A(_01356_ ), .B1(_00636_ ), .B2(_01364_ ), .ZN(_01365_ ) );
INV_X1 _08472_ ( .A(_01298_ ), .ZN(_01366_ ) );
AND2_X1 _08473_ ( .A1(_01366_ ), .A2(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ), .ZN(_01367_ ) );
NOR2_X1 _08474_ ( .A1(_00763_ ), .A2(_01367_ ), .ZN(_01368_ ) );
AND3_X1 _08475_ ( .A1(_00891_ ), .A2(_00785_ ), .A3(\u_exu.acsrd[5] ), .ZN(_01369_ ) );
INV_X1 _08476_ ( .A(_01369_ ), .ZN(_01370_ ) );
INV_X1 _08477_ ( .A(\u_exu.acsrd[8] ), .ZN(_01371_ ) );
NAND3_X1 _08478_ ( .A1(_00785_ ), .A2(_01371_ ), .A3(\u_idu.imm_auipc_lui[28] ), .ZN(_01372_ ) );
NAND3_X1 _08479_ ( .A1(_00862_ ), .A2(_00785_ ), .A3(\u_exu.acsrd[10] ), .ZN(_01373_ ) );
AND3_X1 _08480_ ( .A1(_01370_ ), .A2(_01372_ ), .A3(_01373_ ), .ZN(_01374_ ) );
AOI22_X1 _08481_ ( .A1(_01359_ ), .A2(_00892_ ), .B1(_01355_ ), .B2(_00653_ ), .ZN(_01375_ ) );
AND3_X1 _08482_ ( .A1(_00707_ ), .A2(_00785_ ), .A3(\u_exu.acsrd[7] ), .ZN(_01376_ ) );
AND3_X1 _08483_ ( .A1(_00893_ ), .A2(_00784_ ), .A3(\u_exu.acsrd[3] ), .ZN(_01377_ ) );
INV_X1 _08484_ ( .A(_01377_ ), .ZN(_01378_ ) );
INV_X1 _08485_ ( .A(\u_exu.acsrd[9] ), .ZN(_01379_ ) );
NAND3_X1 _08486_ ( .A1(_00785_ ), .A2(_01379_ ), .A3(\u_idu.imm_auipc_lui[29] ), .ZN(_01380_ ) );
NAND2_X1 _08487_ ( .A1(_01378_ ), .A2(_01380_ ), .ZN(_01381_ ) );
AND2_X1 _08488_ ( .A1(_00785_ ), .A2(\u_exu.acsrd[2] ), .ZN(_01382_ ) );
AOI211_X1 _08489_ ( .A(_01376_ ), .B(_01381_ ), .C1(_00894_ ), .C2(_01382_ ), .ZN(_01383_ ) );
NAND4_X1 _08490_ ( .A1(_01368_ ), .A2(_01374_ ), .A3(_01375_ ), .A4(_01383_ ), .ZN(_01384_ ) );
NOR2_X1 _08491_ ( .A1(ea_err ), .A2(\u_exu.acsrd[6] ), .ZN(_01385_ ) );
INV_X1 _08492_ ( .A(_01385_ ), .ZN(_01386_ ) );
AOI21_X1 _08493_ ( .A(_01386_ ), .B1(_00869_ ), .B2(_00880_ ), .ZN(_01387_ ) );
NOR2_X1 _08494_ ( .A1(_01384_ ), .A2(_01387_ ), .ZN(_01388_ ) );
AND2_X1 _08495_ ( .A1(_01365_ ), .A2(_01388_ ), .ZN(_01389_ ) );
NAND2_X1 _08496_ ( .A1(_00869_ ), .A2(_00880_ ), .ZN(_01390_ ) );
AND2_X1 _08497_ ( .A1(_00636_ ), .A2(_01390_ ), .ZN(_01391_ ) );
NOR2_X1 _08498_ ( .A1(_00633_ ), .A2(\u_idu.imm_auipc_lui[22] ), .ZN(_01392_ ) );
OAI221_X1 _08499_ ( .A(_01389_ ), .B1(_01385_ ), .B2(_01391_ ), .C1(_01382_ ), .C2(_01392_ ), .ZN(_01393_ ) );
AND2_X1 _08500_ ( .A1(_00786_ ), .A2(\u_exu.acsrd[3] ), .ZN(_01394_ ) );
NOR3_X1 _08501_ ( .A1(_00634_ ), .A2(_00893_ ), .A3(_01394_ ), .ZN(_01395_ ) );
INV_X1 _08502_ ( .A(_01395_ ), .ZN(_01396_ ) );
NOR2_X1 _08503_ ( .A1(ea_err ), .A2(\u_exu.acsrd[8] ), .ZN(_01397_ ) );
OR3_X1 _08504_ ( .A1(_00634_ ), .A2(\u_idu.imm_auipc_lui[28] ), .A3(_01397_ ), .ZN(_01398_ ) );
AND2_X1 _08505_ ( .A1(_00785_ ), .A2(\u_exu.acsrd[10] ), .ZN(_01399_ ) );
OR3_X1 _08506_ ( .A1(_00634_ ), .A2(_00862_ ), .A3(_01399_ ), .ZN(_01400_ ) );
NAND3_X1 _08507_ ( .A1(_01396_ ), .A2(_01398_ ), .A3(_01400_ ), .ZN(_01401_ ) );
NOR2_X1 _08508_ ( .A1(_01393_ ), .A2(_01401_ ), .ZN(_01402_ ) );
AND2_X1 _08509_ ( .A1(_00872_ ), .A2(_00635_ ), .ZN(_01403_ ) );
INV_X1 _08510_ ( .A(\u_exu.acsrd[1] ), .ZN(_01404_ ) );
NOR2_X1 _08511_ ( .A1(_01404_ ), .A2(ea_err ), .ZN(_01405_ ) );
XNOR2_X1 _08512_ ( .A(_01403_ ), .B(_01405_ ), .ZN(_01406_ ) );
NAND3_X1 _08513_ ( .A1(_00886_ ), .A2(_00686_ ), .A3(_00713_ ), .ZN(_01407_ ) );
AOI22_X1 _08514_ ( .A1(_01407_ ), .A2(fanout_net_22 ), .B1(_00884_ ), .B2(_00883_ ), .ZN(_01408_ ) );
INV_X1 _08515_ ( .A(_01408_ ), .ZN(_01409_ ) );
NOR2_X1 _08516_ ( .A1(_00634_ ), .A2(_01409_ ), .ZN(_01410_ ) );
NOR2_X1 _08517_ ( .A1(ea_err ), .A2(\u_exu.acsrd[0] ), .ZN(_01411_ ) );
INV_X1 _08518_ ( .A(_01411_ ), .ZN(_01412_ ) );
XNOR2_X1 _08519_ ( .A(_01410_ ), .B(_01412_ ), .ZN(_01413_ ) );
INV_X1 _08520_ ( .A(_01413_ ), .ZN(_01414_ ) );
AND3_X1 _08521_ ( .A1(_01402_ ), .A2(_01406_ ), .A3(_01414_ ), .ZN(_01415_ ) );
BUF_X4 _08522_ ( .A(_01415_ ), .Z(_01416_ ) );
AND2_X1 _08523_ ( .A1(_01113_ ), .A2(_01106_ ), .ZN(_01417_ ) );
NOR2_X2 _08524_ ( .A1(_01417_ ), .A2(_01105_ ), .ZN(_01418_ ) );
NOR2_X2 _08525_ ( .A1(_01418_ ), .A2(_00858_ ), .ZN(_01419_ ) );
INV_X1 _08526_ ( .A(_01419_ ), .ZN(_01420_ ) );
BUF_X4 _08527_ ( .A(_01420_ ), .Z(_01421_ ) );
NAND4_X1 _08528_ ( .A1(_01416_ ), .A2(_00789_ ), .A3(_00788_ ), .A4(_01421_ ), .ZN(_01422_ ) );
NAND3_X1 _08529_ ( .A1(_01402_ ), .A2(_01406_ ), .A3(_01414_ ), .ZN(_01423_ ) );
BUF_X2 _08530_ ( .A(_01423_ ), .Z(_01424_ ) );
BUF_X4 _08531_ ( .A(_01421_ ), .Z(_01425_ ) );
NAND4_X1 _08532_ ( .A1(_00869_ ), .A2(_00880_ ), .A3(_00708_ ), .A4(_00755_ ), .ZN(_01426_ ) );
AND2_X1 _08533_ ( .A1(_00636_ ), .A2(_01426_ ), .ZN(_01427_ ) );
AOI211_X1 _08534_ ( .A(_01392_ ), .B(_01427_ ), .C1(\u_idu.imm_auipc_lui[23] ), .C2(_00636_ ), .ZN(_01428_ ) );
BUF_X4 _08535_ ( .A(_01428_ ), .Z(_01429_ ) );
NOR2_X2 _08536_ ( .A1(_01403_ ), .A2(_01410_ ), .ZN(_01430_ ) );
BUF_X4 _08537_ ( .A(_01430_ ), .Z(_01431_ ) );
NAND3_X1 _08538_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][31] ), .A3(_01431_ ), .ZN(_01432_ ) );
NOR4_X1 _08539_ ( .A1(_00872_ ), .A2(_00858_ ), .A3(\u_idu.imm_auipc_lui[23] ), .A4(\u_idu.imm_auipc_lui[22] ), .ZN(_01433_ ) );
BUF_X2 _08540_ ( .A(_01433_ ), .Z(_01434_ ) );
NOR3_X1 _08541_ ( .A1(_00858_ ), .A2(_01409_ ), .A3(_01426_ ), .ZN(_01435_ ) );
BUF_X2 _08542_ ( .A(_01435_ ), .Z(_01436_ ) );
NAND3_X1 _08543_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][31] ), .A3(_01436_ ), .ZN(_01437_ ) );
AND2_X1 _08544_ ( .A1(_01392_ ), .A2(_00893_ ), .ZN(_01438_ ) );
BUF_X4 _08545_ ( .A(_01438_ ), .Z(_01439_ ) );
BUF_X4 _08546_ ( .A(_01439_ ), .Z(_01440_ ) );
AND4_X1 _08547_ ( .A1(_00708_ ), .A2(_00636_ ), .A3(_00755_ ), .A4(_01390_ ), .ZN(_01441_ ) );
BUF_X4 _08548_ ( .A(_01441_ ), .Z(_01442_ ) );
NAND4_X1 _08549_ ( .A1(_01431_ ), .A2(\u_csr.csr[2][31] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_01443_ ) );
NAND3_X1 _08550_ ( .A1(_01432_ ), .A2(_01437_ ), .A3(_01443_ ), .ZN(_01444_ ) );
NAND3_X1 _08551_ ( .A1(_01424_ ), .A2(_01425_ ), .A3(_01444_ ), .ZN(_01445_ ) );
AOI21_X1 _08552_ ( .A(_01353_ ), .B1(_01422_ ), .B2(_01445_ ), .ZN(_01446_ ) );
NOR2_X1 _08553_ ( .A1(_00741_ ), .A2(_00705_ ), .ZN(_01447_ ) );
AND4_X1 _08554_ ( .A1(_00761_ ), .A2(_01447_ ), .A3(_00739_ ), .A4(_00722_ ), .ZN(_01448_ ) );
AND2_X1 _08555_ ( .A1(_00675_ ), .A2(_01448_ ), .ZN(_01449_ ) );
AND2_X1 _08556_ ( .A1(_01449_ ), .A2(_00747_ ), .ZN(_01450_ ) );
NOR2_X1 _08557_ ( .A1(_01450_ ), .A2(_00743_ ), .ZN(_01451_ ) );
AND3_X1 _08558_ ( .A1(_00675_ ), .A2(_01448_ ), .A3(_00759_ ), .ZN(_01452_ ) );
NOR2_X1 _08559_ ( .A1(_01451_ ), .A2(_01452_ ), .ZN(_01453_ ) );
INV_X1 _08560_ ( .A(_01453_ ), .ZN(_01454_ ) );
BUF_X4 _08561_ ( .A(_01454_ ), .Z(_01455_ ) );
AOI221_X4 _08562_ ( .A(_01446_ ), .B1(\de_pc[31] ), .B2(_01455_ ), .C1(_01063_ ), .C2(_01066_ ), .ZN(_01456_ ) );
AND2_X1 _08563_ ( .A1(_00662_ ), .A2(_00668_ ), .ZN(_01457_ ) );
NOR4_X1 _08564_ ( .A1(_01457_ ), .A2(_00673_ ), .A3(_00734_ ), .A4(_00694_ ), .ZN(_01458_ ) );
AND2_X1 _08565_ ( .A1(_01458_ ), .A2(_01447_ ), .ZN(_01459_ ) );
BUF_X2 _08566_ ( .A(_01459_ ), .Z(_01460_ ) );
OR3_X1 _08567_ ( .A1(_01302_ ), .A2(_01346_ ), .A3(_01460_ ), .ZN(_01461_ ) );
AND2_X1 _08568_ ( .A1(_01459_ ), .A2(_01084_ ), .ZN(_01462_ ) );
BUF_X4 _08569_ ( .A(_01462_ ), .Z(_01463_ ) );
BUF_X4 _08570_ ( .A(_01463_ ), .Z(_01464_ ) );
OAI21_X1 _08571_ ( .A(_00732_ ), .B1(_00665_ ), .B2(_00719_ ), .ZN(_01465_ ) );
AND2_X1 _08572_ ( .A1(_01081_ ), .A2(_01465_ ), .ZN(_01466_ ) );
AND2_X2 _08573_ ( .A1(_01459_ ), .A2(_01466_ ), .ZN(_01467_ ) );
BUF_X4 _08574_ ( .A(_01467_ ), .Z(_01468_ ) );
NOR2_X1 _08575_ ( .A1(_00727_ ), .A2(_00692_ ), .ZN(_01469_ ) );
AND2_X2 _08576_ ( .A1(_01469_ ), .A2(_00924_ ), .ZN(_01470_ ) );
OR2_X1 _08577_ ( .A1(_01470_ ), .A2(_00653_ ), .ZN(_01471_ ) );
AOI21_X1 _08578_ ( .A(_00653_ ), .B1(\u_idu.imm_auipc_lui[12] ), .B2(_00677_ ), .ZN(_01472_ ) );
AND2_X1 _08579_ ( .A1(_00733_ ), .A2(_01472_ ), .ZN(_01473_ ) );
INV_X1 _08580_ ( .A(_01473_ ), .ZN(_01474_ ) );
AND4_X1 _08581_ ( .A1(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A2(_00645_ ), .A3(_00677_ ), .A4(\u_idu.imm_auipc_lui[31] ), .ZN(_01475_ ) );
AND2_X1 _08582_ ( .A1(_00720_ ), .A2(_01475_ ), .ZN(_01476_ ) );
INV_X1 _08583_ ( .A(_01476_ ), .ZN(_01477_ ) );
OAI211_X1 _08584_ ( .A(_00719_ ), .B(\u_idu.imm_auipc_lui[31] ), .C1(_00732_ ), .C2(_00667_ ), .ZN(_01478_ ) );
AND3_X1 _08585_ ( .A1(_01474_ ), .A2(_01477_ ), .A3(_01478_ ), .ZN(_01479_ ) );
NAND2_X1 _08586_ ( .A1(_01471_ ), .A2(_01479_ ), .ZN(_01480_ ) );
AOI221_X4 _08587_ ( .A(_01052_ ), .B1(\de_pc[31] ), .B2(_01464_ ), .C1(_01468_ ), .C2(_01480_ ), .ZN(_01481_ ) );
AOI221_X1 _08588_ ( .A(_00897_ ), .B1(_01347_ ), .B2(_01456_ ), .C1(_01461_ ), .C2(_01481_ ), .ZN(_00129_ ) );
BUF_X4 _08589_ ( .A(_01244_ ), .Z(_01482_ ) );
BUF_X2 _08590_ ( .A(_01320_ ), .Z(_01483_ ) );
BUF_X4 _08591_ ( .A(_00915_ ), .Z(_01484_ ) );
BUF_X4 _08592_ ( .A(_01316_ ), .Z(_01485_ ) );
BUF_X4 _08593_ ( .A(_00909_ ), .Z(_01486_ ) );
AOI22_X1 _08594_ ( .A1(_01485_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01486_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01487_ ) );
BUF_X4 _08595_ ( .A(_01005_ ), .Z(_01488_ ) );
BUF_X4 _08596_ ( .A(_01309_ ), .Z(_01489_ ) );
AOI22_X1 _08597_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01490_ ) );
AOI21_X1 _08598_ ( .A(_01484_ ), .B1(_01487_ ), .B2(_01490_ ), .ZN(_01491_ ) );
BUF_X4 _08599_ ( .A(_01309_ ), .Z(_01492_ ) );
AOI22_X1 _08600_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01493_ ) );
BUF_X4 _08601_ ( .A(_00950_ ), .Z(_01494_ ) );
BUF_X4 _08602_ ( .A(_00909_ ), .Z(_01495_ ) );
AOI22_X1 _08603_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01496_ ) );
AOI21_X1 _08604_ ( .A(_01327_ ), .B1(_01493_ ), .B2(_01496_ ), .ZN(_01497_ ) );
OAI21_X1 _08605_ ( .A(_01483_ ), .B1(_01491_ ), .B2(_01497_ ), .ZN(_01498_ ) );
AOI22_X1 _08606_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01486_ ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01499_ ) );
BUF_X4 _08607_ ( .A(_01337_ ), .Z(_01500_ ) );
NAND3_X1 _08608_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01328_ ), .ZN(_01501_ ) );
NAND3_X1 _08609_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01325_ ), .ZN(_01502_ ) );
NAND4_X1 _08610_ ( .A1(_01499_ ), .A2(_01336_ ), .A3(_01501_ ), .A4(_01502_ ), .ZN(_01503_ ) );
BUF_X2 _08611_ ( .A(_01046_ ), .Z(_01504_ ) );
NAND3_X1 _08612_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01328_ ), .ZN(_01505_ ) );
BUF_X4 _08613_ ( .A(_00976_ ), .Z(_01506_ ) );
INV_X1 _08614_ ( .A(\u_reg.rf[1][30] ), .ZN(_01507_ ) );
AOI21_X1 _08615_ ( .A(_01506_ ), .B1(_01325_ ), .B2(_01507_ ), .ZN(_01508_ ) );
NOR2_X1 _08616_ ( .A1(_01342_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01509_ ) );
OAI211_X1 _08617_ ( .A(_01327_ ), .B(_01505_ ), .C1(_01508_ ), .C2(_01509_ ), .ZN(_01510_ ) );
NAND3_X1 _08618_ ( .A1(_01503_ ), .A2(_01504_ ), .A3(_01510_ ), .ZN(_01511_ ) );
AND2_X1 _08619_ ( .A1(_01498_ ), .A2(_01511_ ), .ZN(_01512_ ) );
OAI21_X1 _08620_ ( .A(_01303_ ), .B1(_01482_ ), .B2(_01512_ ), .ZN(_01513_ ) );
OR2_X1 _08621_ ( .A1(_01212_ ), .A2(\io_master_rdata[30] ), .ZN(_01514_ ) );
INV_X1 _08622_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_31_A_$_ANDNOT__Y_B ), .ZN(_01515_ ) );
OR3_X1 _08623_ ( .A1(_01208_ ), .A2(\u_arbiter.raddr[2] ), .A3(_01515_ ), .ZN(_01516_ ) );
INV_X1 _08624_ ( .A(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .ZN(_01517_ ) );
BUF_X2 _08625_ ( .A(_01208_ ), .Z(_01518_ ) );
OAI21_X1 _08626_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ), .B1(_01518_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_01519_ ) );
NAND3_X1 _08627_ ( .A1(_01516_ ), .A2(_01517_ ), .A3(_01519_ ), .ZN(_01520_ ) );
NAND3_X1 _08628_ ( .A1(_01192_ ), .A2(_01211_ ), .A3(_01520_ ), .ZN(_01521_ ) );
AND2_X1 _08629_ ( .A1(_01514_ ), .A2(_01521_ ), .ZN(_01522_ ) );
BUF_X2 _08630_ ( .A(_01276_ ), .Z(_01523_ ) );
AND3_X1 _08631_ ( .A1(_01522_ ), .A2(_01523_ ), .A3(_01278_ ), .ZN(_01524_ ) );
NOR3_X1 _08632_ ( .A1(_01275_ ), .A2(_01294_ ), .A3(_01524_ ), .ZN(_01525_ ) );
NAND2_X1 _08633_ ( .A1(_01525_ ), .A2(fanout_net_11 ), .ZN(_01526_ ) );
BUF_X4 _08634_ ( .A(_01298_ ), .Z(_01527_ ) );
MUX2_X1 _08635_ ( .A(\ea_addr[30] ), .B(\u_exu.ecsr[30] ), .S(_01527_ ), .Z(_01528_ ) );
OR2_X1 _08636_ ( .A1(_01528_ ), .A2(fanout_net_11 ), .ZN(_01529_ ) );
AND2_X1 _08637_ ( .A1(_01526_ ), .A2(_01529_ ), .ZN(\ar_data[30] ) );
INV_X1 _08638_ ( .A(\ar_data[30] ), .ZN(_01530_ ) );
BUF_X4 _08639_ ( .A(_01304_ ), .Z(_01531_ ) );
AOI21_X1 _08640_ ( .A(_01513_ ), .B1(_01530_ ), .B2(_01531_ ), .ZN(_01532_ ) );
BUF_X2 _08641_ ( .A(_00743_ ), .Z(_01533_ ) );
NAND2_X1 _08642_ ( .A1(_01532_ ), .A2(_01533_ ), .ZN(_01534_ ) );
BUF_X4 _08643_ ( .A(_01352_ ), .Z(_01535_ ) );
NAND4_X1 _08644_ ( .A1(_01416_ ), .A2(_00791_ ), .A3(_00790_ ), .A4(_01421_ ), .ZN(_01536_ ) );
BUF_X4 _08645_ ( .A(_01423_ ), .Z(_01537_ ) );
BUF_X4 _08646_ ( .A(_01420_ ), .Z(_01538_ ) );
AND2_X2 _08647_ ( .A1(_01430_ ), .A2(_01439_ ), .ZN(_01539_ ) );
AND3_X1 _08648_ ( .A1(_00707_ ), .A2(\u_idu.imm_auipc_lui[24] ), .A3(\u_idu.imm_auipc_lui[29] ), .ZN(_01540_ ) );
NAND4_X1 _08649_ ( .A1(_00636_ ), .A2(\u_idu.imm_auipc_lui[31] ), .A3(_00891_ ), .A4(_01540_ ), .ZN(_01541_ ) );
OAI211_X1 _08650_ ( .A(\u_idu.imm_auipc_lui[28] ), .B(\u_idu.imm_auipc_lui[30] ), .C1(_00763_ ), .C2(_00786_ ), .ZN(_01542_ ) );
NOR3_X1 _08651_ ( .A1(_01391_ ), .A2(_01541_ ), .A3(_01542_ ), .ZN(_01543_ ) );
AND2_X2 _08652_ ( .A1(_01539_ ), .A2(_01543_ ), .ZN(_01544_ ) );
INV_X1 _08653_ ( .A(_01544_ ), .ZN(_01545_ ) );
NAND3_X1 _08654_ ( .A1(_01428_ ), .A2(\u_csr.csr[1][30] ), .A3(_01430_ ), .ZN(_01546_ ) );
NOR2_X1 _08655_ ( .A1(_00885_ ), .A2(_00887_ ), .ZN(_01547_ ) );
AOI22_X1 _08656_ ( .A1(_00637_ ), .A2(_01426_ ), .B1(fanout_net_23 ), .B2(_01547_ ), .ZN(_01548_ ) );
NAND4_X1 _08657_ ( .A1(_01440_ ), .A2(\u_csr.csr[0][30] ), .A3(_01410_ ), .A4(_01548_ ), .ZN(_01549_ ) );
NAND4_X1 _08658_ ( .A1(_01430_ ), .A2(\u_csr.csr[2][30] ), .A3(_01439_ ), .A4(_01441_ ), .ZN(_01550_ ) );
NAND4_X1 _08659_ ( .A1(_01545_ ), .A2(_01546_ ), .A3(_01549_ ), .A4(_01550_ ), .ZN(_01551_ ) );
NAND3_X1 _08660_ ( .A1(_01537_ ), .A2(_01538_ ), .A3(_01551_ ), .ZN(_01552_ ) );
AOI21_X1 _08661_ ( .A(_01535_ ), .B1(_01536_ ), .B2(_01552_ ), .ZN(_01553_ ) );
AOI221_X4 _08662_ ( .A(_01553_ ), .B1(\de_pc[30] ), .B2(_01455_ ), .C1(_01063_ ), .C2(_01066_ ), .ZN(_01554_ ) );
INV_X1 _08663_ ( .A(_01460_ ), .ZN(_01555_ ) );
BUF_X4 _08664_ ( .A(_01555_ ), .Z(_01556_ ) );
BUF_X4 _08665_ ( .A(_01556_ ), .Z(_01557_ ) );
NAND2_X1 _08666_ ( .A1(_01532_ ), .A2(_01557_ ), .ZN(_01558_ ) );
OR2_X1 _08667_ ( .A1(_01473_ ), .A2(_01476_ ), .ZN(_01559_ ) );
INV_X1 _08668_ ( .A(_01559_ ), .ZN(_01560_ ) );
AND2_X1 _08669_ ( .A1(_01471_ ), .A2(_01560_ ), .ZN(_01561_ ) );
INV_X1 _08670_ ( .A(_01561_ ), .ZN(_01562_ ) );
BUF_X4 _08671_ ( .A(_00738_ ), .Z(_01563_ ) );
AOI21_X1 _08672_ ( .A(_01562_ ), .B1(\u_idu.imm_auipc_lui[30] ), .B2(_01563_ ), .ZN(_01564_ ) );
INV_X1 _08673_ ( .A(_01466_ ), .ZN(_01565_ ) );
BUF_X4 _08674_ ( .A(_01565_ ), .Z(_01566_ ) );
NOR3_X1 _08675_ ( .A1(_01564_ ), .A2(_01556_ ), .A3(_01566_ ), .ZN(_01567_ ) );
AOI211_X1 _08676_ ( .A(_01567_ ), .B(_01053_ ), .C1(\de_pc[30] ), .C2(_01464_ ), .ZN(_01568_ ) );
AOI221_X4 _08677_ ( .A(_00897_ ), .B1(_01534_ ), .B2(_01554_ ), .C1(_01558_ ), .C2(_01568_ ), .ZN(_00130_ ) );
AOI22_X1 _08678_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01569_ ) );
BUF_X4 _08679_ ( .A(_01005_ ), .Z(_01570_ ) );
AOI22_X1 _08680_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01571_ ) );
NAND3_X1 _08681_ ( .A1(_01569_ ), .A2(_01571_ ), .A3(_01327_ ), .ZN(_01572_ ) );
AOI22_X1 _08682_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01573_ ) );
AOI22_X1 _08683_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01574_ ) );
NAND3_X1 _08684_ ( .A1(_01573_ ), .A2(_01574_ ), .A3(_01318_ ), .ZN(_01575_ ) );
AND3_X1 _08685_ ( .A1(_01572_ ), .A2(_01575_ ), .A3(_01483_ ), .ZN(_01576_ ) );
BUF_X4 _08686_ ( .A(_01323_ ), .Z(_01577_ ) );
OAI211_X1 _08687_ ( .A(fanout_net_21 ), .B(_01322_ ), .C1(_01577_ ), .C2(\u_reg.rf[1][21] ), .ZN(_01578_ ) );
OAI21_X1 _08688_ ( .A(_01578_ ), .B1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01342_ ), .ZN(_01579_ ) );
BUF_X4 _08689_ ( .A(_00975_ ), .Z(_01580_ ) );
NAND4_X1 _08690_ ( .A1(_01328_ ), .A2(fanout_net_21 ), .A3(_01322_ ), .A4(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01581_ ) );
NAND3_X1 _08691_ ( .A1(_01579_ ), .A2(_01580_ ), .A3(_01581_ ), .ZN(_01582_ ) );
AND2_X1 _08692_ ( .A1(_01582_ ), .A2(_01504_ ), .ZN(_01583_ ) );
AOI22_X1 _08693_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01333_ ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01584_ ) );
BUF_X4 _08694_ ( .A(_01484_ ), .Z(_01585_ ) );
BUF_X4 _08695_ ( .A(_01500_ ), .Z(_01586_ ) );
BUF_X4 _08696_ ( .A(_01577_ ), .Z(_01587_ ) );
NAND3_X1 _08697_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01587_ ), .ZN(_01588_ ) );
BUF_X4 _08698_ ( .A(_01341_ ), .Z(_01589_ ) );
NAND3_X1 _08699_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01589_ ), .ZN(_01590_ ) );
NAND4_X1 _08700_ ( .A1(_01584_ ), .A2(_01585_ ), .A3(_01588_ ), .A4(_01590_ ), .ZN(_01591_ ) );
AOI21_X1 _08701_ ( .A(_01576_ ), .B1(_01583_ ), .B2(_01591_ ), .ZN(_01592_ ) );
OAI21_X1 _08702_ ( .A(_01303_ ), .B1(_01482_ ), .B2(_01592_ ), .ZN(_01593_ ) );
OR2_X4 _08703_ ( .A1(_01275_ ), .A2(_01294_ ), .ZN(_01594_ ) );
BUF_X2 _08704_ ( .A(_01278_ ), .Z(\io_master_arsize[1] ) );
BUF_X4 _08705_ ( .A(_01213_ ), .Z(_01595_ ) );
INV_X1 _08706_ ( .A(\u_lsu.u_clint.mtime[21] ), .ZN(_01596_ ) );
NAND4_X1 _08707_ ( .A1(_01276_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_01596_ ), .ZN(_01597_ ) );
BUF_X4 _08708_ ( .A(_01209_ ), .Z(_01598_ ) );
BUF_X4 _08709_ ( .A(_01598_ ), .Z(_01599_ ) );
OAI211_X1 _08710_ ( .A(_01595_ ), .B(_01597_ ), .C1(\u_lsu.u_clint.mtime[53] ), .C2(_01599_ ), .ZN(_01600_ ) );
BUF_X4 _08711_ ( .A(_01214_ ), .Z(_01601_ ) );
NAND2_X1 _08712_ ( .A1(_01601_ ), .A2(\io_master_rdata[21] ), .ZN(_01602_ ) );
AND3_X1 _08713_ ( .A1(_01600_ ), .A2(_01276_ ), .A3(_01602_ ), .ZN(_01603_ ) );
INV_X1 _08714_ ( .A(\u_lsu.u_clint.mtime[29] ), .ZN(_01604_ ) );
NAND4_X1 _08715_ ( .A1(_01252_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_01604_ ), .ZN(_01605_ ) );
OAI211_X1 _08716_ ( .A(_01595_ ), .B(_01605_ ), .C1(\u_lsu.u_clint.mtime[61] ), .C2(_01598_ ), .ZN(_01606_ ) );
NAND2_X1 _08717_ ( .A1(_01214_ ), .A2(\io_master_rdata[29] ), .ZN(_01607_ ) );
AND2_X1 _08718_ ( .A1(_01606_ ), .A2(_01607_ ), .ZN(_01608_ ) );
AOI211_X1 _08719_ ( .A(\io_master_araddr[1] ), .B(_01603_ ), .C1(\io_master_araddr[0] ), .C2(_01608_ ), .ZN(_01609_ ) );
AOI21_X1 _08720_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_01609_ ), .ZN(_01610_ ) );
NAND2_X1 _08721_ ( .A1(_01610_ ), .A2(fanout_net_11 ), .ZN(_01611_ ) );
MUX2_X1 _08722_ ( .A(\ea_addr[21] ), .B(\u_exu.ecsr[21] ), .S(_01527_ ), .Z(_01612_ ) );
OR2_X1 _08723_ ( .A1(_01612_ ), .A2(fanout_net_11 ), .ZN(_01613_ ) );
AND2_X1 _08724_ ( .A1(_01611_ ), .A2(_01613_ ), .ZN(\ar_data[21] ) );
INV_X1 _08725_ ( .A(\ar_data[21] ), .ZN(_01614_ ) );
AOI21_X1 _08726_ ( .A(_01593_ ), .B1(_01614_ ), .B2(_01531_ ), .ZN(_01615_ ) );
NAND2_X1 _08727_ ( .A1(_01615_ ), .A2(_01533_ ), .ZN(_01616_ ) );
AND2_X1 _08728_ ( .A1(_01423_ ), .A2(_01420_ ), .ZN(_01617_ ) );
INV_X1 _08729_ ( .A(_01617_ ), .ZN(_01618_ ) );
BUF_X2 _08730_ ( .A(_01618_ ), .Z(_01619_ ) );
CLKBUF_X2 _08731_ ( .A(_00755_ ), .Z(_01620_ ) );
AND2_X1 _08732_ ( .A1(_01391_ ), .A2(_00708_ ), .ZN(_01621_ ) );
CLKBUF_X2 _08733_ ( .A(_01621_ ), .Z(_01622_ ) );
AND4_X1 _08734_ ( .A1(\u_csr.csr[2][21] ), .A2(_01539_ ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_01623_ ) );
INV_X1 _08735_ ( .A(_01439_ ), .ZN(_01624_ ) );
NAND3_X1 _08736_ ( .A1(_00872_ ), .A2(_00636_ ), .A3(_01408_ ), .ZN(_01625_ ) );
NOR2_X1 _08737_ ( .A1(_01624_ ), .A2(_01625_ ), .ZN(_01626_ ) );
AND2_X2 _08738_ ( .A1(_01626_ ), .A2(_01543_ ), .ZN(_01627_ ) );
NOR3_X1 _08739_ ( .A1(_01623_ ), .A2(_01544_ ), .A3(_01627_ ), .ZN(_01628_ ) );
AND4_X1 _08740_ ( .A1(\u_csr.csr[0][21] ), .A2(_01439_ ), .A3(_01410_ ), .A4(_01548_ ), .ZN(_01629_ ) );
AND2_X1 _08741_ ( .A1(_01428_ ), .A2(_01430_ ), .ZN(_01630_ ) );
BUF_X4 _08742_ ( .A(_01630_ ), .Z(_01631_ ) );
AOI21_X1 _08743_ ( .A(_01629_ ), .B1(_01631_ ), .B2(\u_csr.csr[1][21] ), .ZN(_01632_ ) );
AOI21_X1 _08744_ ( .A(_01619_ ), .B1(_01628_ ), .B2(_01632_ ), .ZN(_01633_ ) );
AOI211_X1 _08745_ ( .A(_01419_ ), .B(_01537_ ), .C1(_00792_ ), .C2(_00793_ ), .ZN(_01634_ ) );
NOR2_X1 _08746_ ( .A1(_01633_ ), .A2(_01634_ ), .ZN(_01635_ ) );
NOR2_X1 _08747_ ( .A1(_01635_ ), .A2(_01353_ ), .ZN(_01636_ ) );
AOI211_X1 _08748_ ( .A(_01077_ ), .B(_01636_ ), .C1(\de_pc[21] ), .C2(_01455_ ), .ZN(_01637_ ) );
NAND2_X1 _08749_ ( .A1(_01615_ ), .A2(_01557_ ), .ZN(_01638_ ) );
BUF_X4 _08750_ ( .A(_00748_ ), .Z(_01639_ ) );
BUF_X4 _08751_ ( .A(_01639_ ), .Z(_01640_ ) );
BUF_X2 _08752_ ( .A(_01640_ ), .Z(_01641_ ) );
OAI21_X1 _08753_ ( .A(_01561_ ), .B1(_01641_ ), .B2(_00928_ ), .ZN(_01642_ ) );
AOI221_X4 _08754_ ( .A(_01052_ ), .B1(\de_pc[21] ), .B2(_01464_ ), .C1(_01468_ ), .C2(_01642_ ), .ZN(_01643_ ) );
AOI221_X1 _08755_ ( .A(_00897_ ), .B1(_01616_ ), .B2(_01637_ ), .C1(_01638_ ), .C2(_01643_ ), .ZN(_00131_ ) );
BUF_X4 _08756_ ( .A(_00896_ ), .Z(_01644_ ) );
AOI22_X1 _08757_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01645_ ) );
AOI22_X1 _08758_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01646_ ) );
NAND3_X1 _08759_ ( .A1(_01645_ ), .A2(_01646_ ), .A3(_01312_ ), .ZN(_01647_ ) );
AOI22_X1 _08760_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01648_ ) );
AOI22_X1 _08761_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01649_ ) );
NAND3_X1 _08762_ ( .A1(_01648_ ), .A2(_01649_ ), .A3(_01318_ ), .ZN(_01650_ ) );
AND3_X1 _08763_ ( .A1(_01647_ ), .A2(_01650_ ), .A3(_01320_ ), .ZN(_01651_ ) );
NAND3_X1 _08764_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01587_ ), .ZN(_01652_ ) );
INV_X1 _08765_ ( .A(\u_reg.rf[1][20] ), .ZN(_01653_ ) );
AOI21_X1 _08766_ ( .A(_01506_ ), .B1(_01589_ ), .B2(_01653_ ), .ZN(_01654_ ) );
NOR2_X1 _08767_ ( .A1(_01589_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01655_ ) );
OAI211_X1 _08768_ ( .A(_01580_ ), .B(_01652_ ), .C1(_01654_ ), .C2(_01655_ ), .ZN(_01656_ ) );
AOI22_X1 _08769_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01486_ ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01657_ ) );
NAND3_X1 _08770_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01577_ ), .ZN(_01658_ ) );
NAND3_X1 _08771_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01325_ ), .ZN(_01659_ ) );
NAND4_X1 _08772_ ( .A1(_01657_ ), .A2(_01484_ ), .A3(_01658_ ), .A4(_01659_ ), .ZN(_01660_ ) );
AND2_X1 _08773_ ( .A1(_01660_ ), .A2(_01504_ ), .ZN(_01661_ ) );
AOI21_X1 _08774_ ( .A(_01651_ ), .B1(_01656_ ), .B2(_01661_ ), .ZN(_01662_ ) );
OAI21_X1 _08775_ ( .A(_01303_ ), .B1(_01482_ ), .B2(_01662_ ), .ZN(_01663_ ) );
BUF_X4 _08776_ ( .A(_01253_ ), .Z(_01664_ ) );
OR2_X1 _08777_ ( .A1(_01212_ ), .A2(\io_master_rdata[20] ), .ZN(_01665_ ) );
BUF_X2 _08778_ ( .A(_01192_ ), .Z(_01666_ ) );
BUF_X2 _08779_ ( .A(_01211_ ), .Z(_01667_ ) );
INV_X1 _08780_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ), .ZN(_01668_ ) );
OR3_X1 _08781_ ( .A1(_01208_ ), .A2(\u_arbiter.raddr[2] ), .A3(_01668_ ), .ZN(_01669_ ) );
BUF_X4 _08782_ ( .A(_01517_ ), .Z(_01670_ ) );
OAI21_X1 _08783_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_10_A_$_ANDNOT__Y_B ), .B1(_01518_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_01671_ ) );
NAND3_X1 _08784_ ( .A1(_01669_ ), .A2(_01670_ ), .A3(_01671_ ), .ZN(_01672_ ) );
NAND3_X1 _08785_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_01672_ ), .ZN(_01673_ ) );
AOI21_X1 _08786_ ( .A(_01664_ ), .B1(_01665_ ), .B2(_01673_ ), .ZN(_01674_ ) );
BUF_X4 _08787_ ( .A(_01664_ ), .Z(_01675_ ) );
INV_X1 _08788_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ), .ZN(_01676_ ) );
OR3_X1 _08789_ ( .A1(_01518_ ), .A2(\u_arbiter.raddr[2] ), .A3(_01676_ ), .ZN(_01677_ ) );
OAI21_X1 _08790_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ), .B1(_01518_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_01678_ ) );
NAND3_X1 _08791_ ( .A1(_01677_ ), .A2(_01670_ ), .A3(_01678_ ), .ZN(_01679_ ) );
NAND3_X1 _08792_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_01679_ ), .ZN(_01680_ ) );
BUF_X2 _08793_ ( .A(_01212_ ), .Z(_01681_ ) );
OAI211_X1 _08794_ ( .A(_01270_ ), .B(_01680_ ), .C1(_01681_ ), .C2(\io_master_rdata[28] ), .ZN(_01682_ ) );
AOI21_X1 _08795_ ( .A(_01674_ ), .B1(_01675_ ), .B2(_01682_ ), .ZN(_01683_ ) );
AOI21_X1 _08796_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_01683_ ), .ZN(_01684_ ) );
NAND2_X1 _08797_ ( .A1(_01684_ ), .A2(fanout_net_11 ), .ZN(_01685_ ) );
MUX2_X1 _08798_ ( .A(\ea_addr[20] ), .B(\u_exu.ecsr[20] ), .S(_01527_ ), .Z(_01686_ ) );
OR2_X1 _08799_ ( .A1(_01686_ ), .A2(fanout_net_11 ), .ZN(_01687_ ) );
AND2_X1 _08800_ ( .A1(_01685_ ), .A2(_01687_ ), .ZN(\ar_data[20] ) );
INV_X1 _08801_ ( .A(\ar_data[20] ), .ZN(_01688_ ) );
AOI21_X1 _08802_ ( .A(_01663_ ), .B1(_01688_ ), .B2(_01531_ ), .ZN(_01689_ ) );
NAND2_X1 _08803_ ( .A1(_01689_ ), .A2(_01533_ ), .ZN(_01690_ ) );
AND3_X1 _08804_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][20] ), .A3(_01435_ ), .ZN(_01691_ ) );
INV_X1 _08805_ ( .A(_01627_ ), .ZN(_01692_ ) );
NAND4_X1 _08806_ ( .A1(_01539_ ), .A2(\u_csr.csr[2][20] ), .A3(_00755_ ), .A4(_01621_ ), .ZN(_01693_ ) );
NAND3_X1 _08807_ ( .A1(_01545_ ), .A2(_01692_ ), .A3(_01693_ ), .ZN(_01694_ ) );
AOI211_X1 _08808_ ( .A(_01691_ ), .B(_01694_ ), .C1(\u_csr.csr[1][20] ), .C2(_01630_ ), .ZN(_01695_ ) );
OR2_X1 _08809_ ( .A1(_01618_ ), .A2(_01695_ ), .ZN(_01696_ ) );
INV_X1 _08810_ ( .A(_01382_ ), .ZN(_01697_ ) );
XNOR2_X1 _08811_ ( .A(_01392_ ), .B(_01697_ ), .ZN(_01698_ ) );
AND3_X1 _08812_ ( .A1(_01698_ ), .A2(_01396_ ), .A3(_01378_ ), .ZN(_01699_ ) );
NAND3_X1 _08813_ ( .A1(_01406_ ), .A2(_01699_ ), .A3(_01414_ ), .ZN(_01700_ ) );
OR3_X1 _08814_ ( .A1(_00634_ ), .A2(\u_idu.imm_auipc_lui[29] ), .A3(_01363_ ), .ZN(_01701_ ) );
AND4_X1 _08815_ ( .A1(_01398_ ), .A2(_01701_ ), .A3(_01372_ ), .A4(_01380_ ), .ZN(_01702_ ) );
AOI21_X1 _08816_ ( .A(_01356_ ), .B1(_00653_ ), .B2(_01355_ ), .ZN(_01703_ ) );
NAND4_X1 _08817_ ( .A1(_01702_ ), .A2(_01703_ ), .A3(_01400_ ), .A4(_01373_ ), .ZN(_01704_ ) );
AOI21_X1 _08818_ ( .A(_01385_ ), .B1(_00636_ ), .B2(_01390_ ), .ZN(_01705_ ) );
NOR3_X1 _08819_ ( .A1(_00634_ ), .A2(_00707_ ), .A3(_01362_ ), .ZN(_01706_ ) );
NOR4_X1 _08820_ ( .A1(_01705_ ), .A2(_01706_ ), .A3(_01387_ ), .A4(_01376_ ), .ZN(_01707_ ) );
NOR2_X1 _08821_ ( .A1(_00634_ ), .A2(_00892_ ), .ZN(_01708_ ) );
XNOR2_X1 _08822_ ( .A(_01708_ ), .B(_01359_ ), .ZN(_01709_ ) );
NAND3_X1 _08823_ ( .A1(_00636_ ), .A2(\u_idu.imm_auipc_lui[25] ), .A3(_01358_ ), .ZN(_01710_ ) );
NAND4_X1 _08824_ ( .A1(_01707_ ), .A2(_01370_ ), .A3(_01709_ ), .A4(_01710_ ), .ZN(_01711_ ) );
NOR3_X1 _08825_ ( .A1(_01700_ ), .A2(_01704_ ), .A3(_01711_ ), .ZN(_01712_ ) );
AND2_X1 _08826_ ( .A1(_01712_ ), .A2(_01368_ ), .ZN(_01713_ ) );
NAND4_X1 _08827_ ( .A1(_01713_ ), .A2(_00795_ ), .A3(_00794_ ), .A4(_01421_ ), .ZN(_01714_ ) );
AOI21_X1 _08828_ ( .A(_01535_ ), .B1(_01696_ ), .B2(_01714_ ), .ZN(_01715_ ) );
AOI221_X4 _08829_ ( .A(_01715_ ), .B1(\de_pc[20] ), .B2(_01455_ ), .C1(_01066_ ), .C2(_01062_ ), .ZN(_01716_ ) );
NAND2_X1 _08830_ ( .A1(_01689_ ), .A2(_01557_ ), .ZN(_01717_ ) );
OAI21_X1 _08831_ ( .A(_01561_ ), .B1(_00878_ ), .B2(_00928_ ), .ZN(_01718_ ) );
AOI221_X4 _08832_ ( .A(_01052_ ), .B1(\de_pc[20] ), .B2(_01463_ ), .C1(_01468_ ), .C2(_01718_ ), .ZN(_01719_ ) );
AOI221_X1 _08833_ ( .A(_01644_ ), .B1(_01690_ ), .B2(_01716_ ), .C1(_01717_ ), .C2(_01719_ ), .ZN(_00132_ ) );
NOR2_X1 _08834_ ( .A1(_01077_ ), .A2(_00896_ ), .ZN(_01720_ ) );
BUF_X4 _08835_ ( .A(_01720_ ), .Z(_01721_ ) );
AND3_X1 _08836_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[19] ), .ZN(_01722_ ) );
BUF_X4 _08837_ ( .A(_01366_ ), .Z(_01723_ ) );
AOI211_X1 _08838_ ( .A(fanout_net_11 ), .B(_01722_ ), .C1(_01723_ ), .C2(\ea_addr[19] ), .ZN(_01724_ ) );
INV_X1 _08839_ ( .A(\u_lsu.u_clint.mtime[19] ), .ZN(_01725_ ) );
NAND4_X1 _08840_ ( .A1(_01276_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_01725_ ), .ZN(_01726_ ) );
OAI211_X1 _08841_ ( .A(_01595_ ), .B(_01726_ ), .C1(\u_lsu.u_clint.mtime[51] ), .C2(_01599_ ), .ZN(_01727_ ) );
NAND2_X1 _08842_ ( .A1(_01601_ ), .A2(\io_master_rdata[19] ), .ZN(_01728_ ) );
AND3_X1 _08843_ ( .A1(_01727_ ), .A2(_01523_ ), .A3(_01728_ ), .ZN(_01729_ ) );
INV_X1 _08844_ ( .A(\u_lsu.u_clint.mtime[27] ), .ZN(_01730_ ) );
NAND4_X1 _08845_ ( .A1(_01276_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_01730_ ), .ZN(_01731_ ) );
OAI211_X1 _08846_ ( .A(_01595_ ), .B(_01731_ ), .C1(\u_lsu.u_clint.mtime[59] ), .C2(_01599_ ), .ZN(_01732_ ) );
NAND2_X1 _08847_ ( .A1(_01601_ ), .A2(\io_master_rdata[27] ), .ZN(_01733_ ) );
AND2_X1 _08848_ ( .A1(_01732_ ), .A2(_01733_ ), .ZN(_01734_ ) );
AOI211_X1 _08849_ ( .A(\io_master_araddr[1] ), .B(_01729_ ), .C1(\io_master_araddr[0] ), .C2(_01734_ ), .ZN(_01735_ ) );
AOI21_X1 _08850_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_01735_ ), .ZN(_01736_ ) );
AOI21_X1 _08851_ ( .A(_01724_ ), .B1(_01736_ ), .B2(fanout_net_11 ), .ZN(\ar_data[19] ) );
NOR2_X1 _08852_ ( .A1(\ar_data[19] ), .A2(_01246_ ), .ZN(_01737_ ) );
BUF_X4 _08853_ ( .A(_01485_ ), .Z(_01738_ ) );
BUF_X4 _08854_ ( .A(_01486_ ), .Z(_01739_ ) );
AOI22_X1 _08855_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01740_ ) );
BUF_X4 _08856_ ( .A(_01488_ ), .Z(_01741_ ) );
BUF_X4 _08857_ ( .A(_01489_ ), .Z(_01742_ ) );
AOI22_X1 _08858_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01743_ ) );
BUF_X2 _08859_ ( .A(_01484_ ), .Z(_01744_ ) );
NAND3_X1 _08860_ ( .A1(_01740_ ), .A2(_01743_ ), .A3(_01744_ ), .ZN(_01745_ ) );
BUF_X2 _08861_ ( .A(_01327_ ), .Z(_01746_ ) );
BUF_X4 _08862_ ( .A(_01338_ ), .Z(_01747_ ) );
BUF_X4 _08863_ ( .A(_01339_ ), .Z(_01748_ ) );
NAND3_X1 _08864_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01748_ ), .ZN(_01749_ ) );
BUF_X4 _08865_ ( .A(_01342_ ), .Z(_01750_ ) );
INV_X1 _08866_ ( .A(\u_reg.rf[1][19] ), .ZN(_01751_ ) );
AOI21_X1 _08867_ ( .A(_01506_ ), .B1(_01750_ ), .B2(_01751_ ), .ZN(_01752_ ) );
NOR2_X1 _08868_ ( .A1(_01750_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01753_ ) );
OAI211_X1 _08869_ ( .A(_01746_ ), .B(_01749_ ), .C1(_01752_ ), .C2(_01753_ ), .ZN(_01754_ ) );
NAND3_X1 _08870_ ( .A1(_01745_ ), .A2(_01504_ ), .A3(_01754_ ), .ZN(_01755_ ) );
BUF_X2 _08871_ ( .A(_01483_ ), .Z(_01756_ ) );
BUF_X4 _08872_ ( .A(_01485_ ), .Z(_01757_ ) );
BUF_X4 _08873_ ( .A(_01486_ ), .Z(_01758_ ) );
AOI22_X1 _08874_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01759_ ) );
BUF_X4 _08875_ ( .A(_01570_ ), .Z(_01760_ ) );
BUF_X4 _08876_ ( .A(_01489_ ), .Z(_01761_ ) );
AOI22_X1 _08877_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01762_ ) );
AOI21_X1 _08878_ ( .A(_01585_ ), .B1(_01759_ ), .B2(_01762_ ), .ZN(_01763_ ) );
AOI22_X1 _08879_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01764_ ) );
AOI22_X1 _08880_ ( .A1(_01485_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01333_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01765_ ) );
AOI21_X1 _08881_ ( .A(_01746_ ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_01766_ ) );
OAI21_X1 _08882_ ( .A(_01756_ ), .B1(_01763_ ), .B2(_01766_ ), .ZN(_01767_ ) );
AOI21_X1 _08883_ ( .A(_01482_ ), .B1(_01755_ ), .B2(_01767_ ), .ZN(_01768_ ) );
OR3_X1 _08884_ ( .A1(_01737_ ), .A2(_00735_ ), .A3(_01768_ ), .ZN(_01769_ ) );
BUF_X4 _08885_ ( .A(_00723_ ), .Z(_01770_ ) );
NOR2_X1 _08886_ ( .A1(_01769_ ), .A2(_01770_ ), .ZN(_01771_ ) );
BUF_X2 _08887_ ( .A(_01416_ ), .Z(_01772_ ) );
BUF_X4 _08888_ ( .A(_01425_ ), .Z(_01773_ ) );
NAND4_X1 _08889_ ( .A1(_01772_ ), .A2(_00799_ ), .A3(_00798_ ), .A4(_01773_ ), .ZN(_01774_ ) );
NAND2_X1 _08890_ ( .A1(_01712_ ), .A2(_01368_ ), .ZN(_01775_ ) );
BUF_X2 _08891_ ( .A(_01775_ ), .Z(_01776_ ) );
BUF_X2 _08892_ ( .A(_01425_ ), .Z(_01777_ ) );
BUF_X4 _08893_ ( .A(_01428_ ), .Z(_01778_ ) );
BUF_X4 _08894_ ( .A(_01430_ ), .Z(_01779_ ) );
BUF_X4 _08895_ ( .A(_01779_ ), .Z(_01780_ ) );
NAND3_X1 _08896_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][19] ), .A3(_01780_ ), .ZN(_01781_ ) );
AND3_X1 _08897_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][19] ), .A3(_01436_ ), .ZN(_01782_ ) );
BUF_X4 _08898_ ( .A(_01543_ ), .Z(_01783_ ) );
AOI21_X1 _08899_ ( .A(_01782_ ), .B1(_01783_ ), .B2(_01626_ ), .ZN(_01784_ ) );
BUF_X4 _08900_ ( .A(_01439_ ), .Z(_01785_ ) );
BUF_X4 _08901_ ( .A(_01441_ ), .Z(_01786_ ) );
NAND4_X1 _08902_ ( .A1(_01780_ ), .A2(\u_csr.csr[2][19] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_01787_ ) );
NAND3_X1 _08903_ ( .A1(_01781_ ), .A2(_01784_ ), .A3(_01787_ ), .ZN(_01788_ ) );
NAND3_X1 _08904_ ( .A1(_01776_ ), .A2(_01777_ ), .A3(_01788_ ), .ZN(_01789_ ) );
AND2_X1 _08905_ ( .A1(_01774_ ), .A2(_01789_ ), .ZN(_01790_ ) );
BUF_X4 _08906_ ( .A(_01353_ ), .Z(_01791_ ) );
INV_X1 _08907_ ( .A(\de_pc[19] ), .ZN(_01792_ ) );
BUF_X4 _08908_ ( .A(_01453_ ), .Z(_01793_ ) );
OAI22_X1 _08909_ ( .A1(_01790_ ), .A2(_01791_ ), .B1(_01792_ ), .B2(_01793_ ), .ZN(_01794_ ) );
OAI21_X1 _08910_ ( .A(_01721_ ), .B1(_01771_ ), .B2(_01794_ ), .ZN(_01795_ ) );
BUF_X4 _08911_ ( .A(_01460_ ), .Z(_01796_ ) );
INV_X2 _08912_ ( .A(_01464_ ), .ZN(_01797_ ) );
OAI22_X1 _08913_ ( .A1(_01769_ ), .A2(_01796_ ), .B1(_01792_ ), .B2(_01797_ ), .ZN(_01798_ ) );
OAI21_X1 _08914_ ( .A(\u_idu.imm_auipc_lui[19] ), .B1(_00746_ ), .B2(_01563_ ), .ZN(_01799_ ) );
OAI21_X1 _08915_ ( .A(\u_idu.imm_auipc_lui[31] ), .B1(_00726_ ), .B2(_00692_ ), .ZN(_01800_ ) );
AND3_X1 _08916_ ( .A1(_01560_ ), .A2(_01799_ ), .A3(_01800_ ), .ZN(_01801_ ) );
INV_X1 _08917_ ( .A(_01801_ ), .ZN(_01802_ ) );
AOI21_X1 _08918_ ( .A(_01798_ ), .B1(_01468_ ), .B2(_01802_ ), .ZN(_01803_ ) );
AND2_X1 _08919_ ( .A1(_01050_ ), .A2(_00895_ ), .ZN(_01804_ ) );
INV_X1 _08920_ ( .A(_01804_ ), .ZN(_01805_ ) );
BUF_X4 _08921_ ( .A(_01805_ ), .Z(_01806_ ) );
OAI21_X1 _08922_ ( .A(_01795_ ), .B1(_01803_ ), .B2(_01806_ ), .ZN(_00133_ ) );
BUF_X2 _08923_ ( .A(_01804_ ), .Z(_00302_ ) );
AND3_X1 _08924_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[18] ), .ZN(_01807_ ) );
AOI211_X1 _08925_ ( .A(fanout_net_11 ), .B(_01807_ ), .C1(_01723_ ), .C2(\ea_addr[18] ), .ZN(_01808_ ) );
OR2_X1 _08926_ ( .A1(_01212_ ), .A2(\io_master_rdata[18] ), .ZN(_01809_ ) );
NAND2_X1 _08927_ ( .A1(_01598_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ), .ZN(_01810_ ) );
OAI21_X1 _08928_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ), .B1(_01208_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_01811_ ) );
NAND3_X1 _08929_ ( .A1(_01810_ ), .A2(_01517_ ), .A3(_01811_ ), .ZN(_01812_ ) );
NAND3_X1 _08930_ ( .A1(_01192_ ), .A2(_01211_ ), .A3(_01812_ ), .ZN(_01813_ ) );
AND2_X1 _08931_ ( .A1(_01809_ ), .A2(_01813_ ), .ZN(_01814_ ) );
OR2_X1 _08932_ ( .A1(_01212_ ), .A2(\io_master_rdata[26] ), .ZN(_01815_ ) );
NAND2_X1 _08933_ ( .A1(_01209_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ), .ZN(_01816_ ) );
OAI21_X1 _08934_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ), .B1(_01208_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_01817_ ) );
NAND3_X1 _08935_ ( .A1(_01816_ ), .A2(_01517_ ), .A3(_01817_ ), .ZN(_01818_ ) );
NAND3_X1 _08936_ ( .A1(_01192_ ), .A2(_01211_ ), .A3(_01818_ ), .ZN(_01819_ ) );
AND3_X1 _08937_ ( .A1(_01815_ ), .A2(_01270_ ), .A3(_01819_ ), .ZN(_01820_ ) );
MUX2_X1 _08938_ ( .A(_01814_ ), .B(_01820_ ), .S(_01675_ ), .Z(_01821_ ) );
AOI21_X1 _08939_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_01821_ ), .ZN(_01822_ ) );
AOI21_X1 _08940_ ( .A(_01808_ ), .B1(_01822_ ), .B2(fanout_net_11 ), .ZN(\ar_data[18] ) );
BUF_X2 _08941_ ( .A(_01245_ ), .Z(_01823_ ) );
OR2_X1 _08942_ ( .A1(\ar_data[18] ), .A2(_01823_ ), .ZN(_01824_ ) );
BUF_X4 _08943_ ( .A(_01246_ ), .Z(_01825_ ) );
BUF_X4 _08944_ ( .A(_01758_ ), .Z(_01826_ ) );
BUF_X4 _08945_ ( .A(_01761_ ), .Z(_01827_ ) );
AOI22_X1 _08946_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01826_ ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01828_ ) );
BUF_X2 _08947_ ( .A(_01585_ ), .Z(_01829_ ) );
BUF_X4 _08948_ ( .A(_01586_ ), .Z(_01830_ ) );
BUF_X4 _08949_ ( .A(_01587_ ), .Z(_01831_ ) );
NAND3_X1 _08950_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_01832_ ) );
BUF_X4 _08951_ ( .A(_01589_ ), .Z(_01833_ ) );
NAND3_X1 _08952_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01833_ ), .ZN(_01834_ ) );
NAND4_X1 _08953_ ( .A1(_01828_ ), .A2(_01829_ ), .A3(_01832_ ), .A4(_01834_ ), .ZN(_01835_ ) );
BUF_X2 _08954_ ( .A(_01504_ ), .Z(_01836_ ) );
BUF_X4 _08955_ ( .A(_00902_ ), .Z(_01837_ ) );
BUF_X4 _08956_ ( .A(_01837_ ), .Z(_01838_ ) );
OAI211_X1 _08957_ ( .A(fanout_net_21 ), .B(_01838_ ), .C1(_01748_ ), .C2(\u_reg.rf[1][18] ), .ZN(_01839_ ) );
OAI21_X1 _08958_ ( .A(_01839_ ), .B1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01833_ ), .ZN(_01840_ ) );
BUF_X2 _08959_ ( .A(_01580_ ), .Z(_01841_ ) );
NAND4_X1 _08960_ ( .A1(_01831_ ), .A2(fanout_net_21 ), .A3(_01838_ ), .A4(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01842_ ) );
NAND3_X1 _08961_ ( .A1(_01840_ ), .A2(_01841_ ), .A3(_01842_ ), .ZN(_01843_ ) );
AND3_X1 _08962_ ( .A1(_01835_ ), .A2(_01836_ ), .A3(_01843_ ), .ZN(_01844_ ) );
BUF_X4 _08963_ ( .A(_01485_ ), .Z(_01845_ ) );
AOI22_X1 _08964_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01826_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01846_ ) );
BUF_X4 _08965_ ( .A(_01760_ ), .Z(_01847_ ) );
AOI22_X1 _08966_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01848_ ) );
NAND3_X1 _08967_ ( .A1(_01846_ ), .A2(_01848_ ), .A3(_01841_ ), .ZN(_01849_ ) );
BUF_X4 _08968_ ( .A(_01334_ ), .Z(_01850_ ) );
AOI22_X1 _08969_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01851_ ) );
BUF_X4 _08970_ ( .A(_01333_ ), .Z(_01852_ ) );
AOI22_X1 _08971_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01853_ ) );
NAND3_X1 _08972_ ( .A1(_01851_ ), .A2(_01853_ ), .A3(_01829_ ), .ZN(_01854_ ) );
BUF_X2 _08973_ ( .A(_01483_ ), .Z(_01855_ ) );
AND3_X1 _08974_ ( .A1(_01849_ ), .A2(_01854_ ), .A3(_01855_ ), .ZN(_01856_ ) );
OAI21_X1 _08975_ ( .A(_01825_ ), .B1(_01844_ ), .B2(_01856_ ), .ZN(_01857_ ) );
NAND3_X1 _08976_ ( .A1(_01824_ ), .A2(_01303_ ), .A3(_01857_ ), .ZN(_01858_ ) );
INV_X1 _08977_ ( .A(\de_pc[18] ), .ZN(_01859_ ) );
OAI22_X1 _08978_ ( .A1(_01858_ ), .A2(_01796_ ), .B1(_01859_ ), .B2(_01797_ ), .ZN(_01860_ ) );
BUF_X2 _08979_ ( .A(_01566_ ), .Z(_01861_ ) );
AND2_X1 _08980_ ( .A1(_01560_ ), .A2(_01800_ ), .ZN(_01862_ ) );
INV_X1 _08981_ ( .A(_01862_ ), .ZN(_01863_ ) );
NOR2_X1 _08982_ ( .A1(_00746_ ), .A2(_01563_ ), .ZN(_01864_ ) );
INV_X1 _08983_ ( .A(_01864_ ), .ZN(_01865_ ) );
AOI21_X1 _08984_ ( .A(_01863_ ), .B1(\u_idu.imm_auipc_lui[18] ), .B2(_01865_ ), .ZN(_01866_ ) );
NOR3_X1 _08985_ ( .A1(_01557_ ), .A2(_01861_ ), .A3(_01866_ ), .ZN(_01867_ ) );
OAI21_X1 _08986_ ( .A(_00302_ ), .B1(_01860_ ), .B2(_01867_ ), .ZN(_01868_ ) );
BUF_X4 _08987_ ( .A(_01720_ ), .Z(_01869_ ) );
NOR2_X1 _08988_ ( .A1(_01858_ ), .A2(_01770_ ), .ZN(_01870_ ) );
NAND4_X1 _08989_ ( .A1(_01772_ ), .A2(_00801_ ), .A3(_00800_ ), .A4(_01777_ ), .ZN(_01871_ ) );
NAND3_X1 _08990_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][18] ), .A3(_01779_ ), .ZN(_01872_ ) );
BUF_X2 _08991_ ( .A(_01434_ ), .Z(_01873_ ) );
BUF_X2 _08992_ ( .A(_01436_ ), .Z(_01874_ ) );
NAND3_X1 _08993_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][18] ), .A3(_01874_ ), .ZN(_01875_ ) );
NAND4_X1 _08994_ ( .A1(_01779_ ), .A2(\u_csr.csr[2][18] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_01876_ ) );
NAND4_X1 _08995_ ( .A1(_01692_ ), .A2(_01872_ ), .A3(_01875_ ), .A4(_01876_ ), .ZN(_01877_ ) );
NAND3_X1 _08996_ ( .A1(_01424_ ), .A2(_01777_ ), .A3(_01877_ ), .ZN(_01878_ ) );
AND2_X1 _08997_ ( .A1(_01871_ ), .A2(_01878_ ), .ZN(_01879_ ) );
OAI22_X1 _08998_ ( .A1(_01879_ ), .A2(_01791_ ), .B1(_01859_ ), .B2(_01793_ ), .ZN(_01880_ ) );
OAI21_X1 _08999_ ( .A(_01869_ ), .B1(_01870_ ), .B2(_01880_ ), .ZN(_01881_ ) );
NAND2_X1 _09000_ ( .A1(_01868_ ), .A2(_01881_ ), .ZN(_00134_ ) );
AND3_X1 _09001_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[17] ), .ZN(_01882_ ) );
AOI211_X1 _09002_ ( .A(fanout_net_11 ), .B(_01882_ ), .C1(_01723_ ), .C2(\ea_addr[17] ), .ZN(_01883_ ) );
BUF_X4 _09003_ ( .A(_01285_ ), .Z(_01884_ ) );
INV_X1 _09004_ ( .A(\u_lsu.u_clint.mtime[25] ), .ZN(_01885_ ) );
NAND4_X1 _09005_ ( .A1(_01276_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_01885_ ), .ZN(_01886_ ) );
OAI211_X1 _09006_ ( .A(_01595_ ), .B(_01886_ ), .C1(\u_lsu.u_clint.mtime[57] ), .C2(_01599_ ), .ZN(_01887_ ) );
NAND2_X1 _09007_ ( .A1(_01601_ ), .A2(\io_master_rdata[25] ), .ZN(_01888_ ) );
AOI21_X1 _09008_ ( .A(_01884_ ), .B1(_01887_ ), .B2(_01888_ ), .ZN(_01889_ ) );
INV_X1 _09009_ ( .A(\u_lsu.u_clint.mtime[17] ), .ZN(_01890_ ) );
NAND4_X1 _09010_ ( .A1(_01276_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_01890_ ), .ZN(_01891_ ) );
OAI211_X1 _09011_ ( .A(_01595_ ), .B(_01891_ ), .C1(\u_lsu.u_clint.mtime[49] ), .C2(_01598_ ), .ZN(_01892_ ) );
NAND2_X1 _09012_ ( .A1(_01601_ ), .A2(\io_master_rdata[17] ), .ZN(_01893_ ) );
AND2_X1 _09013_ ( .A1(_01892_ ), .A2(_01893_ ), .ZN(_01894_ ) );
INV_X1 _09014_ ( .A(_01894_ ), .ZN(_01895_ ) );
MUX2_X1 _09015_ ( .A(_01889_ ), .B(_01895_ ), .S(_01523_ ), .Z(_01896_ ) );
AOI21_X1 _09016_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_01896_ ), .ZN(_01897_ ) );
AOI21_X1 _09017_ ( .A(_01883_ ), .B1(_01897_ ), .B2(fanout_net_11 ), .ZN(\ar_data[17] ) );
OR2_X1 _09018_ ( .A1(\ar_data[17] ), .A2(_01823_ ), .ZN(_01898_ ) );
BUF_X4 _09019_ ( .A(_01334_ ), .Z(_01899_ ) );
AOI22_X1 _09020_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01852_ ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01900_ ) );
BUF_X4 _09021_ ( .A(_01336_ ), .Z(_01901_ ) );
BUF_X4 _09022_ ( .A(_01338_ ), .Z(_01902_ ) );
BUF_X4 _09023_ ( .A(_01339_ ), .Z(_01903_ ) );
NAND3_X1 _09024_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01903_ ), .ZN(_01904_ ) );
BUF_X4 _09025_ ( .A(_01342_ ), .Z(_01905_ ) );
NAND3_X1 _09026_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01905_ ), .ZN(_01906_ ) );
NAND4_X1 _09027_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(_01904_ ), .A4(_01906_ ), .ZN(_01907_ ) );
OAI211_X1 _09028_ ( .A(fanout_net_21 ), .B(_01838_ ), .C1(_01748_ ), .C2(\u_reg.rf[1][17] ), .ZN(_01908_ ) );
OAI21_X1 _09029_ ( .A(_01908_ ), .B1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01833_ ), .ZN(_01909_ ) );
BUF_X2 _09030_ ( .A(_01580_ ), .Z(_01910_ ) );
NAND4_X1 _09031_ ( .A1(_01831_ ), .A2(fanout_net_21 ), .A3(_01838_ ), .A4(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01911_ ) );
NAND3_X1 _09032_ ( .A1(_01909_ ), .A2(_01910_ ), .A3(_01911_ ), .ZN(_01912_ ) );
AND3_X1 _09033_ ( .A1(_01907_ ), .A2(_01836_ ), .A3(_01912_ ), .ZN(_01913_ ) );
BUF_X4 _09034_ ( .A(_01485_ ), .Z(_01914_ ) );
BUF_X4 _09035_ ( .A(_01333_ ), .Z(_01915_ ) );
AOI22_X1 _09036_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01915_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01916_ ) );
BUF_X4 _09037_ ( .A(_01488_ ), .Z(_01917_ ) );
AOI22_X1 _09038_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01918_ ) );
NAND3_X1 _09039_ ( .A1(_01916_ ), .A2(_01918_ ), .A3(_01901_ ), .ZN(_01919_ ) );
AOI22_X1 _09040_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01920_ ) );
AOI22_X1 _09041_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01921_ ) );
NAND3_X1 _09042_ ( .A1(_01920_ ), .A2(_01921_ ), .A3(_01910_ ), .ZN(_01922_ ) );
AND3_X1 _09043_ ( .A1(_01919_ ), .A2(_01922_ ), .A3(_01855_ ), .ZN(_01923_ ) );
OAI21_X1 _09044_ ( .A(_01823_ ), .B1(_01913_ ), .B2(_01923_ ), .ZN(_01924_ ) );
NAND3_X1 _09045_ ( .A1(_01898_ ), .A2(_01303_ ), .A3(_01924_ ), .ZN(_01925_ ) );
NOR2_X1 _09046_ ( .A1(_01925_ ), .A2(_01770_ ), .ZN(_01926_ ) );
AND3_X1 _09047_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][17] ), .A3(_01436_ ), .ZN(_01927_ ) );
BUF_X2 _09048_ ( .A(_01539_ ), .Z(_01928_ ) );
NAND4_X1 _09049_ ( .A1(_01928_ ), .A2(\u_csr.csr[2][17] ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_01929_ ) );
NAND3_X1 _09050_ ( .A1(_01545_ ), .A2(_01692_ ), .A3(_01929_ ), .ZN(_01930_ ) );
AOI211_X1 _09051_ ( .A(_01927_ ), .B(_01930_ ), .C1(\u_csr.csr[1][17] ), .C2(_01631_ ), .ZN(_01931_ ) );
OR2_X1 _09052_ ( .A1(_01619_ ), .A2(_01931_ ), .ZN(_01932_ ) );
NAND4_X1 _09053_ ( .A1(_01713_ ), .A2(_00803_ ), .A3(_00802_ ), .A4(_01773_ ), .ZN(_01933_ ) );
AND2_X1 _09054_ ( .A1(_01932_ ), .A2(_01933_ ), .ZN(_01934_ ) );
INV_X1 _09055_ ( .A(\de_pc[17] ), .ZN(_01935_ ) );
OAI22_X1 _09056_ ( .A1(_01934_ ), .A2(_01791_ ), .B1(_01935_ ), .B2(_01793_ ), .ZN(_01936_ ) );
OAI21_X1 _09057_ ( .A(_01721_ ), .B1(_01926_ ), .B2(_01936_ ), .ZN(_01937_ ) );
OAI22_X1 _09058_ ( .A1(_01925_ ), .A2(_01796_ ), .B1(_01935_ ), .B2(_01797_ ), .ZN(_01938_ ) );
OAI21_X1 _09059_ ( .A(\u_idu.imm_auipc_lui[17] ), .B1(_00746_ ), .B2(_01563_ ), .ZN(_01939_ ) );
AND3_X1 _09060_ ( .A1(_01560_ ), .A2(_01800_ ), .A3(_01939_ ), .ZN(_01940_ ) );
INV_X1 _09061_ ( .A(_01940_ ), .ZN(_01941_ ) );
AOI21_X1 _09062_ ( .A(_01938_ ), .B1(_01468_ ), .B2(_01941_ ), .ZN(_01942_ ) );
OAI21_X1 _09063_ ( .A(_01937_ ), .B1(_01942_ ), .B2(_01806_ ), .ZN(_00135_ ) );
AND3_X1 _09064_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[16] ), .ZN(_01943_ ) );
AOI211_X1 _09065_ ( .A(fanout_net_11 ), .B(_01943_ ), .C1(_01723_ ), .C2(\ea_addr[16] ), .ZN(_01944_ ) );
OR2_X1 _09066_ ( .A1(_01681_ ), .A2(\io_master_rdata[16] ), .ZN(_01945_ ) );
BUF_X2 _09067_ ( .A(_01518_ ), .Z(_01946_ ) );
INV_X1 _09068_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ), .ZN(_01947_ ) );
OR3_X1 _09069_ ( .A1(_01946_ ), .A2(\u_arbiter.raddr[2] ), .A3(_01947_ ), .ZN(_01948_ ) );
OAI21_X1 _09070_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ), .B1(_01946_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_01949_ ) );
NAND3_X1 _09071_ ( .A1(_01948_ ), .A2(_01670_ ), .A3(_01949_ ), .ZN(_01950_ ) );
NAND3_X1 _09072_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_01950_ ), .ZN(_01951_ ) );
AOI21_X1 _09073_ ( .A(_01664_ ), .B1(_01945_ ), .B2(_01951_ ), .ZN(_01952_ ) );
OR2_X1 _09074_ ( .A1(_01681_ ), .A2(\io_master_rdata[24] ), .ZN(_01953_ ) );
INV_X1 _09075_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ), .ZN(_01954_ ) );
OR3_X1 _09076_ ( .A1(_01518_ ), .A2(\u_arbiter.raddr[2] ), .A3(_01954_ ), .ZN(_01955_ ) );
OAI21_X1 _09077_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ), .B1(_01946_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_01956_ ) );
NAND3_X1 _09078_ ( .A1(_01955_ ), .A2(_01670_ ), .A3(_01956_ ), .ZN(_01957_ ) );
NAND3_X1 _09079_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_01957_ ), .ZN(_01958_ ) );
AND2_X1 _09080_ ( .A1(_01953_ ), .A2(_01958_ ), .ZN(_01959_ ) );
INV_X1 _09081_ ( .A(_01959_ ), .ZN(_01960_ ) );
AOI211_X1 _09082_ ( .A(\io_master_araddr[1] ), .B(_01952_ ), .C1(_01960_ ), .C2(\io_master_araddr[0] ), .ZN(_01961_ ) );
AOI21_X1 _09083_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_01961_ ), .ZN(_01962_ ) );
AOI21_X1 _09084_ ( .A(_01944_ ), .B1(_01962_ ), .B2(fanout_net_11 ), .ZN(\ar_data[16] ) );
NOR2_X1 _09085_ ( .A1(\ar_data[16] ), .A2(_01246_ ), .ZN(_01963_ ) );
AOI22_X1 _09086_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01739_ ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01964_ ) );
NAND3_X1 _09087_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01748_ ), .ZN(_01965_ ) );
NAND3_X1 _09088_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01750_ ), .ZN(_01966_ ) );
NAND4_X1 _09089_ ( .A1(_01964_ ), .A2(_01744_ ), .A3(_01965_ ), .A4(_01966_ ), .ZN(_01967_ ) );
OAI211_X1 _09090_ ( .A(fanout_net_21 ), .B(_01837_ ), .C1(_01339_ ), .C2(\u_reg.rf[1][16] ), .ZN(_01968_ ) );
OAI21_X1 _09091_ ( .A(_01968_ ), .B1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01750_ ), .ZN(_01969_ ) );
NAND4_X1 _09092_ ( .A1(_01748_ ), .A2(fanout_net_21 ), .A3(_01838_ ), .A4(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01970_ ) );
NAND3_X1 _09093_ ( .A1(_01969_ ), .A2(_01746_ ), .A3(_01970_ ), .ZN(_01971_ ) );
NAND3_X1 _09094_ ( .A1(_01967_ ), .A2(_01504_ ), .A3(_01971_ ), .ZN(_01972_ ) );
AOI22_X1 _09095_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01973_ ) );
AOI22_X1 _09096_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01974_ ) );
AOI21_X1 _09097_ ( .A(_01585_ ), .B1(_01973_ ), .B2(_01974_ ), .ZN(_01975_ ) );
AOI22_X1 _09098_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01976_ ) );
AOI22_X1 _09099_ ( .A1(_01485_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01333_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01977_ ) );
AOI21_X1 _09100_ ( .A(_01580_ ), .B1(_01976_ ), .B2(_01977_ ), .ZN(_01978_ ) );
OAI21_X1 _09101_ ( .A(_01756_ ), .B1(_01975_ ), .B2(_01978_ ), .ZN(_01979_ ) );
AOI21_X1 _09102_ ( .A(_01482_ ), .B1(_01972_ ), .B2(_01979_ ), .ZN(_01980_ ) );
OR3_X1 _09103_ ( .A1(_01963_ ), .A2(_00735_ ), .A3(_01980_ ), .ZN(_01981_ ) );
NOR2_X1 _09104_ ( .A1(_01981_ ), .A2(_01770_ ), .ZN(_01982_ ) );
NAND4_X1 _09105_ ( .A1(_01772_ ), .A2(_00805_ ), .A3(_00804_ ), .A4(_01773_ ), .ZN(_01983_ ) );
AND3_X1 _09106_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][16] ), .A3(_01874_ ), .ZN(_01984_ ) );
AOI21_X1 _09107_ ( .A(_01984_ ), .B1(_01928_ ), .B2(_01783_ ), .ZN(_01985_ ) );
NAND3_X1 _09108_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][16] ), .A3(_01780_ ), .ZN(_01986_ ) );
NAND4_X1 _09109_ ( .A1(_01780_ ), .A2(\u_csr.csr[2][16] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_01987_ ) );
NAND3_X1 _09110_ ( .A1(_01985_ ), .A2(_01986_ ), .A3(_01987_ ), .ZN(_01988_ ) );
NAND3_X1 _09111_ ( .A1(_01776_ ), .A2(_01777_ ), .A3(_01988_ ), .ZN(_01989_ ) );
AND2_X1 _09112_ ( .A1(_01983_ ), .A2(_01989_ ), .ZN(_01990_ ) );
INV_X1 _09113_ ( .A(\de_pc[16] ), .ZN(_01991_ ) );
OAI22_X1 _09114_ ( .A1(_01990_ ), .A2(_01791_ ), .B1(_01991_ ), .B2(_01793_ ), .ZN(_01992_ ) );
OAI21_X1 _09115_ ( .A(_01721_ ), .B1(_01982_ ), .B2(_01992_ ), .ZN(_01993_ ) );
OAI22_X1 _09116_ ( .A1(_01981_ ), .A2(_01796_ ), .B1(_01991_ ), .B2(_01797_ ), .ZN(_01994_ ) );
OAI21_X1 _09117_ ( .A(\u_idu.imm_auipc_lui[16] ), .B1(_00746_ ), .B2(_01563_ ), .ZN(_01995_ ) );
AND3_X1 _09118_ ( .A1(_01560_ ), .A2(_01800_ ), .A3(_01995_ ), .ZN(_01996_ ) );
INV_X1 _09119_ ( .A(_01996_ ), .ZN(_01997_ ) );
AOI21_X1 _09120_ ( .A(_01994_ ), .B1(_01468_ ), .B2(_01997_ ), .ZN(_01998_ ) );
OAI21_X1 _09121_ ( .A(_01993_ ), .B1(_01998_ ), .B2(_01806_ ), .ZN(_00136_ ) );
BUF_X2 _09122_ ( .A(_00735_ ), .Z(_01999_ ) );
AOI22_X1 _09123_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02000_ ) );
AOI22_X1 _09124_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02001_ ) );
NAND3_X1 _09125_ ( .A1(_02000_ ), .A2(_02001_ ), .A3(_01910_ ), .ZN(_02002_ ) );
AOI22_X1 _09126_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02003_ ) );
AOI22_X1 _09127_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01915_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02004_ ) );
NAND3_X1 _09128_ ( .A1(_02003_ ), .A2(_02004_ ), .A3(_01901_ ), .ZN(_02005_ ) );
NAND3_X1 _09129_ ( .A1(_02002_ ), .A2(_02005_ ), .A3(_01855_ ), .ZN(_02006_ ) );
AOI22_X1 _09130_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01915_ ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02007_ ) );
NAND3_X1 _09131_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01903_ ), .ZN(_02008_ ) );
NAND3_X1 _09132_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01905_ ), .ZN(_02009_ ) );
NAND4_X1 _09133_ ( .A1(_02007_ ), .A2(_01901_ ), .A3(_02008_ ), .A4(_02009_ ), .ZN(_02010_ ) );
OAI211_X1 _09134_ ( .A(fanout_net_21 ), .B(_01837_ ), .C1(_01587_ ), .C2(\u_reg.rf[1][15] ), .ZN(_02011_ ) );
OAI21_X1 _09135_ ( .A(_02011_ ), .B1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01905_ ), .ZN(_02012_ ) );
INV_X1 _09136_ ( .A(_01494_ ), .ZN(_02013_ ) );
INV_X1 _09137_ ( .A(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02014_ ) );
OAI211_X1 _09138_ ( .A(_01910_ ), .B(_02012_ ), .C1(_02013_ ), .C2(_02014_ ), .ZN(_02015_ ) );
NAND3_X1 _09139_ ( .A1(_02010_ ), .A2(_01836_ ), .A3(_02015_ ), .ZN(_02016_ ) );
NAND2_X1 _09140_ ( .A1(_02006_ ), .A2(_02016_ ), .ZN(_02017_ ) );
AOI21_X1 _09141_ ( .A(_01999_ ), .B1(_01825_ ), .B2(_02017_ ), .ZN(_02018_ ) );
AND3_X1 _09142_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[15] ), .ZN(_02019_ ) );
AOI211_X1 _09143_ ( .A(fanout_net_11 ), .B(_02019_ ), .C1(_01723_ ), .C2(\ea_addr[15] ), .ZN(_02020_ ) );
AOI21_X1 _09144_ ( .A(_01277_ ), .B1(_01254_ ), .B2(_01271_ ), .ZN(_02021_ ) );
NOR2_X1 _09145_ ( .A1(_01295_ ), .A2(_02021_ ), .ZN(_02022_ ) );
AOI21_X1 _09146_ ( .A(_02020_ ), .B1(_02022_ ), .B2(fanout_net_11 ), .ZN(\ar_data[15] ) );
OAI21_X1 _09147_ ( .A(_02018_ ), .B1(\ar_data[15] ), .B2(_01825_ ), .ZN(_02023_ ) );
NOR2_X1 _09148_ ( .A1(_02023_ ), .A2(_01770_ ), .ZN(_02024_ ) );
NAND4_X1 _09149_ ( .A1(_01772_ ), .A2(_00808_ ), .A3(_00806_ ), .A4(_01773_ ), .ZN(_02025_ ) );
NAND3_X1 _09150_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][15] ), .A3(_01780_ ), .ZN(_02026_ ) );
NAND3_X1 _09151_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][15] ), .A3(_01874_ ), .ZN(_02027_ ) );
NAND4_X1 _09152_ ( .A1(_01780_ ), .A2(\u_csr.csr[2][15] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_02028_ ) );
NAND3_X1 _09153_ ( .A1(_02026_ ), .A2(_02027_ ), .A3(_02028_ ), .ZN(_02029_ ) );
NAND3_X1 _09154_ ( .A1(_01424_ ), .A2(_01777_ ), .A3(_02029_ ), .ZN(_02030_ ) );
AND2_X1 _09155_ ( .A1(_02025_ ), .A2(_02030_ ), .ZN(_02031_ ) );
INV_X1 _09156_ ( .A(\de_pc[15] ), .ZN(_02032_ ) );
OAI22_X1 _09157_ ( .A1(_02031_ ), .A2(_01791_ ), .B1(_02032_ ), .B2(_01793_ ), .ZN(_02033_ ) );
OAI21_X1 _09158_ ( .A(_01721_ ), .B1(_02024_ ), .B2(_02033_ ), .ZN(_02034_ ) );
OAI22_X1 _09159_ ( .A1(_02023_ ), .A2(_01796_ ), .B1(_02032_ ), .B2(_01797_ ), .ZN(_02035_ ) );
OAI21_X1 _09160_ ( .A(fanout_net_21 ), .B1(_00746_ ), .B2(_01563_ ), .ZN(_02036_ ) );
AND3_X1 _09161_ ( .A1(_01560_ ), .A2(_01800_ ), .A3(_02036_ ), .ZN(_02037_ ) );
INV_X1 _09162_ ( .A(_02037_ ), .ZN(_02038_ ) );
AOI21_X1 _09163_ ( .A(_02035_ ), .B1(_01468_ ), .B2(_02038_ ), .ZN(_02039_ ) );
OAI21_X1 _09164_ ( .A(_02034_ ), .B1(_02039_ ), .B2(_01806_ ), .ZN(_00137_ ) );
AOI22_X1 _09165_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01915_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02040_ ) );
AOI22_X1 _09166_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02041_ ) );
NAND3_X1 _09167_ ( .A1(_02040_ ), .A2(_02041_ ), .A3(_01910_ ), .ZN(_02042_ ) );
AOI22_X1 _09168_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02043_ ) );
AOI22_X1 _09169_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02044_ ) );
NAND3_X1 _09170_ ( .A1(_02043_ ), .A2(_02044_ ), .A3(_01901_ ), .ZN(_02045_ ) );
NAND3_X1 _09171_ ( .A1(_02042_ ), .A2(_02045_ ), .A3(_01756_ ), .ZN(_02046_ ) );
AOI22_X1 _09172_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01486_ ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02047_ ) );
NAND3_X1 _09173_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01339_ ), .ZN(_02048_ ) );
NAND3_X1 _09174_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01342_ ), .ZN(_02049_ ) );
AND4_X1 _09175_ ( .A1(_01336_ ), .A2(_02047_ ), .A3(_02048_ ), .A4(_02049_ ), .ZN(_02050_ ) );
OR2_X1 _09176_ ( .A1(_02050_ ), .A2(_01756_ ), .ZN(_02051_ ) );
OR2_X1 _09177_ ( .A1(_01325_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02052_ ) );
OAI211_X1 _09178_ ( .A(fanout_net_21 ), .B(_01837_ ), .C1(_01328_ ), .C2(\u_reg.rf[1][14] ), .ZN(_02053_ ) );
AOI221_X4 _09179_ ( .A(_01336_ ), .B1(_02052_ ), .B2(_02053_ ), .C1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_01757_ ), .ZN(_02054_ ) );
OAI21_X1 _09180_ ( .A(_02046_ ), .B1(_02051_ ), .B2(_02054_ ), .ZN(_02055_ ) );
AOI21_X1 _09181_ ( .A(_01999_ ), .B1(_01825_ ), .B2(_02055_ ), .ZN(_02056_ ) );
AND3_X1 _09182_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[14] ), .ZN(_02057_ ) );
AOI211_X1 _09183_ ( .A(fanout_net_11 ), .B(_02057_ ), .C1(_01723_ ), .C2(\ea_addr[14] ), .ZN(_02058_ ) );
INV_X1 _09184_ ( .A(_01277_ ), .ZN(_02059_ ) );
AND3_X1 _09185_ ( .A1(_01514_ ), .A2(_01255_ ), .A3(_01521_ ), .ZN(_02060_ ) );
OR2_X1 _09186_ ( .A1(_01212_ ), .A2(\io_master_rdata[22] ), .ZN(_02061_ ) );
INV_X1 _09187_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_39_A_$_ANDNOT__Y_B ), .ZN(_02062_ ) );
OR3_X1 _09188_ ( .A1(_01208_ ), .A2(\u_arbiter.raddr[2] ), .A3(_02062_ ), .ZN(_02063_ ) );
OAI21_X1 _09189_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_8_A_$_ANDNOT__Y_B ), .B1(_01518_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_02064_ ) );
NAND3_X1 _09190_ ( .A1(_02063_ ), .A2(_01670_ ), .A3(_02064_ ), .ZN(_02065_ ) );
NAND3_X1 _09191_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_02065_ ), .ZN(_02066_ ) );
AND2_X1 _09192_ ( .A1(_02061_ ), .A2(_02066_ ), .ZN(_02067_ ) );
AOI21_X1 _09193_ ( .A(_02060_ ), .B1(_01270_ ), .B2(_02067_ ), .ZN(_02068_ ) );
NAND2_X1 _09194_ ( .A1(_01599_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ), .ZN(_02069_ ) );
OAI21_X1 _09195_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ), .B1(_01946_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_02070_ ) );
NAND3_X1 _09196_ ( .A1(_02069_ ), .A2(_01670_ ), .A3(_02070_ ), .ZN(_02071_ ) );
NAND3_X1 _09197_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_02071_ ), .ZN(_02072_ ) );
OAI21_X1 _09198_ ( .A(_02072_ ), .B1(_01681_ ), .B2(\io_master_rdata[14] ), .ZN(_02073_ ) );
OAI21_X1 _09199_ ( .A(_02068_ ), .B1(_01675_ ), .B2(_02073_ ), .ZN(_02074_ ) );
AOI21_X1 _09200_ ( .A(_01295_ ), .B1(_02059_ ), .B2(_02074_ ), .ZN(_02075_ ) );
AOI21_X1 _09201_ ( .A(_02058_ ), .B1(_02075_ ), .B2(fanout_net_11 ), .ZN(\ar_data[14] ) );
OAI21_X1 _09202_ ( .A(_02056_ ), .B1(\ar_data[14] ), .B2(_01825_ ), .ZN(_02076_ ) );
NOR2_X1 _09203_ ( .A1(_02076_ ), .A2(_01770_ ), .ZN(_02077_ ) );
NAND4_X1 _09204_ ( .A1(_01772_ ), .A2(_00810_ ), .A3(_00809_ ), .A4(_01773_ ), .ZN(_02078_ ) );
AND3_X1 _09205_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][14] ), .A3(_01874_ ), .ZN(_02079_ ) );
AOI21_X1 _09206_ ( .A(_02079_ ), .B1(_01928_ ), .B2(_01783_ ), .ZN(_02080_ ) );
NAND3_X1 _09207_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][14] ), .A3(_01780_ ), .ZN(_02081_ ) );
NAND4_X1 _09208_ ( .A1(_01779_ ), .A2(\u_csr.csr[2][14] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_02082_ ) );
NAND3_X1 _09209_ ( .A1(_02080_ ), .A2(_02081_ ), .A3(_02082_ ), .ZN(_02083_ ) );
NAND3_X1 _09210_ ( .A1(_01776_ ), .A2(_01777_ ), .A3(_02083_ ), .ZN(_02084_ ) );
AND2_X1 _09211_ ( .A1(_02078_ ), .A2(_02084_ ), .ZN(_02085_ ) );
INV_X1 _09212_ ( .A(\de_pc[14] ), .ZN(_02086_ ) );
OAI22_X1 _09213_ ( .A1(_02085_ ), .A2(_01791_ ), .B1(_02086_ ), .B2(_01793_ ), .ZN(_02087_ ) );
OAI21_X1 _09214_ ( .A(_01721_ ), .B1(_02077_ ), .B2(_02087_ ), .ZN(_02088_ ) );
OAI22_X1 _09215_ ( .A1(_02076_ ), .A2(_01796_ ), .B1(_02086_ ), .B2(_01797_ ), .ZN(_02089_ ) );
AOI21_X1 _09216_ ( .A(_01863_ ), .B1(\u_idu.imm_auipc_lui[14] ), .B2(_01865_ ), .ZN(_02090_ ) );
INV_X1 _09217_ ( .A(_02090_ ), .ZN(_02091_ ) );
AOI21_X1 _09218_ ( .A(_02089_ ), .B1(_01468_ ), .B2(_02091_ ), .ZN(_02092_ ) );
OAI21_X1 _09219_ ( .A(_02088_ ), .B1(_02092_ ), .B2(_01806_ ), .ZN(_00138_ ) );
AOI22_X1 _09220_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02093_ ) );
AOI22_X1 _09221_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02094_ ) );
AOI21_X1 _09222_ ( .A(_01744_ ), .B1(_02093_ ), .B2(_02094_ ), .ZN(_02095_ ) );
AOI22_X1 _09223_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02096_ ) );
AOI22_X1 _09224_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02097_ ) );
AOI21_X1 _09225_ ( .A(_01746_ ), .B1(_02096_ ), .B2(_02097_ ), .ZN(_02098_ ) );
OAI21_X1 _09226_ ( .A(_01756_ ), .B1(_02095_ ), .B2(_02098_ ), .ZN(_02099_ ) );
OR2_X1 _09227_ ( .A1(_01325_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02100_ ) );
OAI211_X1 _09228_ ( .A(fanout_net_21 ), .B(_01837_ ), .C1(_01328_ ), .C2(\u_reg.rf[1][13] ), .ZN(_02101_ ) );
AOI221_X4 _09229_ ( .A(_01336_ ), .B1(_02100_ ), .B2(_02101_ ), .C1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_01738_ ), .ZN(_02102_ ) );
AOI22_X1 _09230_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01915_ ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02103_ ) );
NAND3_X1 _09231_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01903_ ), .ZN(_02104_ ) );
NAND3_X1 _09232_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01905_ ), .ZN(_02105_ ) );
NAND4_X1 _09233_ ( .A1(_02103_ ), .A2(_01744_ ), .A3(_02104_ ), .A4(_02105_ ), .ZN(_02106_ ) );
NAND2_X1 _09234_ ( .A1(_02106_ ), .A2(_01836_ ), .ZN(_02107_ ) );
OAI21_X1 _09235_ ( .A(_02099_ ), .B1(_02102_ ), .B2(_02107_ ), .ZN(_02108_ ) );
AOI21_X1 _09236_ ( .A(_01999_ ), .B1(_01825_ ), .B2(_02108_ ), .ZN(_02109_ ) );
AND3_X1 _09237_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[13] ), .ZN(_02110_ ) );
AOI211_X1 _09238_ ( .A(fanout_net_11 ), .B(_02110_ ), .C1(_01723_ ), .C2(\ea_addr[13] ), .ZN(_02111_ ) );
AOI21_X1 _09239_ ( .A(_01884_ ), .B1(_01600_ ), .B2(_01602_ ), .ZN(_02112_ ) );
AOI21_X1 _09240_ ( .A(_01256_ ), .B1(_01606_ ), .B2(_01607_ ), .ZN(_02113_ ) );
NOR3_X1 _09241_ ( .A1(_01518_ ), .A2(\u_arbiter.raddr[2] ), .A3(\u_lsu.u_clint.mtime[13] ), .ZN(_02114_ ) );
INV_X1 _09242_ ( .A(\u_lsu.u_clint.mtime[45] ), .ZN(_02115_ ) );
INV_X1 _09243_ ( .A(_01598_ ), .ZN(_02116_ ) );
AOI211_X1 _09244_ ( .A(_02114_ ), .B(_01248_ ), .C1(_02115_ ), .C2(_02116_ ), .ZN(_02117_ ) );
AOI21_X1 _09245_ ( .A(_02117_ ), .B1(_01601_ ), .B2(\io_master_rdata[13] ), .ZN(_02118_ ) );
NOR2_X1 _09246_ ( .A1(_02118_ ), .A2(_01675_ ), .ZN(_02119_ ) );
OR3_X1 _09247_ ( .A1(_02112_ ), .A2(_02113_ ), .A3(_02119_ ), .ZN(_02120_ ) );
AOI21_X1 _09248_ ( .A(_01295_ ), .B1(_02059_ ), .B2(_02120_ ), .ZN(_02121_ ) );
AOI21_X1 _09249_ ( .A(_02111_ ), .B1(_02121_ ), .B2(fanout_net_11 ), .ZN(\ar_data[13] ) );
OAI21_X1 _09250_ ( .A(_02109_ ), .B1(\ar_data[13] ), .B2(_01825_ ), .ZN(_02122_ ) );
NOR2_X1 _09251_ ( .A1(_02122_ ), .A2(_01770_ ), .ZN(_02123_ ) );
NAND4_X1 _09252_ ( .A1(_01772_ ), .A2(_00812_ ), .A3(_00811_ ), .A4(_01773_ ), .ZN(_02124_ ) );
AND3_X1 _09253_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][13] ), .A3(_01874_ ), .ZN(_02125_ ) );
AOI21_X1 _09254_ ( .A(_02125_ ), .B1(_01928_ ), .B2(_01783_ ), .ZN(_02126_ ) );
NAND3_X1 _09255_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][13] ), .A3(_01780_ ), .ZN(_02127_ ) );
NAND4_X1 _09256_ ( .A1(_01779_ ), .A2(\u_csr.csr[2][13] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_02128_ ) );
NAND3_X1 _09257_ ( .A1(_02126_ ), .A2(_02127_ ), .A3(_02128_ ), .ZN(_02129_ ) );
NAND3_X1 _09258_ ( .A1(_01776_ ), .A2(_01777_ ), .A3(_02129_ ), .ZN(_02130_ ) );
AND2_X1 _09259_ ( .A1(_02124_ ), .A2(_02130_ ), .ZN(_02131_ ) );
INV_X1 _09260_ ( .A(\de_pc[13] ), .ZN(_02132_ ) );
OAI22_X1 _09261_ ( .A1(_02131_ ), .A2(_01791_ ), .B1(_02132_ ), .B2(_01793_ ), .ZN(_02133_ ) );
OAI21_X1 _09262_ ( .A(_01721_ ), .B1(_02123_ ), .B2(_02133_ ), .ZN(_02134_ ) );
OAI22_X1 _09263_ ( .A1(_02122_ ), .A2(_01796_ ), .B1(_02132_ ), .B2(_01797_ ), .ZN(_02135_ ) );
AOI21_X1 _09264_ ( .A(_01863_ ), .B1(\u_idu.imm_auipc_lui[13] ), .B2(_01865_ ), .ZN(_02136_ ) );
INV_X1 _09265_ ( .A(_02136_ ), .ZN(_02137_ ) );
AOI21_X1 _09266_ ( .A(_02135_ ), .B1(_01468_ ), .B2(_02137_ ), .ZN(_02138_ ) );
OAI21_X1 _09267_ ( .A(_02134_ ), .B1(_02138_ ), .B2(_01806_ ), .ZN(_00139_ ) );
AOI22_X1 _09268_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01915_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02139_ ) );
AOI22_X1 _09269_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02140_ ) );
AOI21_X1 _09270_ ( .A(_01901_ ), .B1(_02139_ ), .B2(_02140_ ), .ZN(_02141_ ) );
AOI22_X1 _09271_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02142_ ) );
AOI22_X1 _09272_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01915_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02143_ ) );
AOI21_X1 _09273_ ( .A(_01910_ ), .B1(_02142_ ), .B2(_02143_ ), .ZN(_02144_ ) );
OAI21_X1 _09274_ ( .A(_01855_ ), .B1(_02141_ ), .B2(_02144_ ), .ZN(_02145_ ) );
AOI22_X1 _09275_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02146_ ) );
AOI22_X1 _09276_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02147_ ) );
AOI21_X1 _09277_ ( .A(_01746_ ), .B1(_02146_ ), .B2(_02147_ ), .ZN(_02148_ ) );
OAI211_X1 _09278_ ( .A(fanout_net_21 ), .B(_01838_ ), .C1(_01748_ ), .C2(\u_reg.rf[1][12] ), .ZN(_02149_ ) );
OAI21_X1 _09279_ ( .A(_02149_ ), .B1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01905_ ), .ZN(_02150_ ) );
INV_X1 _09280_ ( .A(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02151_ ) );
OAI21_X1 _09281_ ( .A(_02150_ ), .B1(_02013_ ), .B2(_02151_ ), .ZN(_02152_ ) );
AOI21_X1 _09282_ ( .A(_02148_ ), .B1(_01841_ ), .B2(_02152_ ), .ZN(_02153_ ) );
OAI21_X1 _09283_ ( .A(_02145_ ), .B1(_02153_ ), .B2(_01855_ ), .ZN(_02154_ ) );
AOI21_X1 _09284_ ( .A(_01999_ ), .B1(_01825_ ), .B2(_02154_ ), .ZN(_02155_ ) );
AND3_X1 _09285_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[12] ), .ZN(_02156_ ) );
AOI211_X1 _09286_ ( .A(fanout_net_11 ), .B(_02156_ ), .C1(_01723_ ), .C2(\ea_addr[12] ), .ZN(_02157_ ) );
AND3_X1 _09287_ ( .A1(_01665_ ), .A2(_01270_ ), .A3(_01673_ ), .ZN(_02158_ ) );
OR2_X1 _09288_ ( .A1(_01681_ ), .A2(\io_master_rdata[28] ), .ZN(_02159_ ) );
AND2_X1 _09289_ ( .A1(_02159_ ), .A2(_01680_ ), .ZN(_02160_ ) );
AOI21_X1 _09290_ ( .A(_02158_ ), .B1(_01255_ ), .B2(_02160_ ), .ZN(_02161_ ) );
NAND2_X1 _09291_ ( .A1(_01598_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ), .ZN(_02162_ ) );
OAI21_X1 _09292_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_18_A_$_ANDNOT__Y_B ), .B1(_01946_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_02163_ ) );
NAND3_X1 _09293_ ( .A1(_02162_ ), .A2(_01670_ ), .A3(_02163_ ), .ZN(_02164_ ) );
NAND3_X1 _09294_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_02164_ ), .ZN(_02165_ ) );
OAI21_X1 _09295_ ( .A(_02165_ ), .B1(_01681_ ), .B2(\io_master_rdata[12] ), .ZN(_02166_ ) );
OAI21_X1 _09296_ ( .A(_02161_ ), .B1(_01675_ ), .B2(_02166_ ), .ZN(_02167_ ) );
AOI21_X1 _09297_ ( .A(_01295_ ), .B1(_02059_ ), .B2(_02167_ ), .ZN(_02168_ ) );
AOI21_X1 _09298_ ( .A(_02157_ ), .B1(_02168_ ), .B2(fanout_net_11 ), .ZN(\ar_data[12] ) );
OAI21_X1 _09299_ ( .A(_02155_ ), .B1(\ar_data[12] ), .B2(_01825_ ), .ZN(_02169_ ) );
INV_X1 _09300_ ( .A(\de_pc[12] ), .ZN(_02170_ ) );
OAI22_X1 _09301_ ( .A1(_02169_ ), .A2(_01796_ ), .B1(_02170_ ), .B2(_01797_ ), .ZN(_02171_ ) );
AOI21_X1 _09302_ ( .A(_01863_ ), .B1(\u_idu.imm_auipc_lui[12] ), .B2(_01865_ ), .ZN(_02172_ ) );
NOR3_X1 _09303_ ( .A1(_01557_ ), .A2(_01861_ ), .A3(_02172_ ), .ZN(_02173_ ) );
OAI21_X1 _09304_ ( .A(_00302_ ), .B1(_02171_ ), .B2(_02173_ ), .ZN(_02174_ ) );
NOR2_X1 _09305_ ( .A1(_02169_ ), .A2(_01770_ ), .ZN(_02175_ ) );
AND3_X1 _09306_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][12] ), .A3(_01436_ ), .ZN(_02176_ ) );
NAND4_X1 _09307_ ( .A1(_01928_ ), .A2(\u_csr.csr[2][12] ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_02177_ ) );
NAND3_X1 _09308_ ( .A1(_01545_ ), .A2(_01692_ ), .A3(_02177_ ), .ZN(_02178_ ) );
AOI211_X1 _09309_ ( .A(_02176_ ), .B(_02178_ ), .C1(\u_csr.csr[1][12] ), .C2(_01631_ ), .ZN(_02179_ ) );
NOR2_X1 _09310_ ( .A1(_01619_ ), .A2(_02179_ ), .ZN(_02180_ ) );
AOI211_X1 _09311_ ( .A(_01419_ ), .B(_01776_ ), .C1(_00852_ ), .C2(_00853_ ), .ZN(_02181_ ) );
NOR2_X1 _09312_ ( .A1(_02180_ ), .A2(_02181_ ), .ZN(_02182_ ) );
OAI22_X1 _09313_ ( .A1(_02182_ ), .A2(_01791_ ), .B1(_02170_ ), .B2(_01793_ ), .ZN(_02183_ ) );
OAI21_X1 _09314_ ( .A(_01869_ ), .B1(_02175_ ), .B2(_02183_ ), .ZN(_02184_ ) );
NAND2_X1 _09315_ ( .A1(_02174_ ), .A2(_02184_ ), .ZN(_00140_ ) );
AOI21_X1 _09316_ ( .A(_01279_ ), .B1(_01606_ ), .B2(_01607_ ), .ZN(_02185_ ) );
NOR3_X1 _09317_ ( .A1(_01275_ ), .A2(_01295_ ), .A3(_02185_ ), .ZN(_02186_ ) );
NAND2_X1 _09318_ ( .A1(_02186_ ), .A2(fanout_net_11 ), .ZN(_02187_ ) );
MUX2_X1 _09319_ ( .A(\ea_addr[29] ), .B(\u_exu.ecsr[29] ), .S(_01299_ ), .Z(_02188_ ) );
OR2_X1 _09320_ ( .A1(_02188_ ), .A2(fanout_net_12 ), .ZN(_02189_ ) );
AOI21_X1 _09321_ ( .A(_01246_ ), .B1(_02187_ ), .B2(_02189_ ), .ZN(_02190_ ) );
AOI22_X1 _09322_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02191_ ) );
AOI22_X1 _09323_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02192_ ) );
NAND3_X1 _09324_ ( .A1(_02191_ ), .A2(_02192_ ), .A3(_01312_ ), .ZN(_02193_ ) );
AOI22_X1 _09325_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02194_ ) );
AOI22_X1 _09326_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02195_ ) );
NAND3_X1 _09327_ ( .A1(_02194_ ), .A2(_02195_ ), .A3(_01318_ ), .ZN(_02196_ ) );
AND3_X1 _09328_ ( .A1(_02193_ ), .A2(_02196_ ), .A3(_01320_ ), .ZN(_02197_ ) );
OAI211_X1 _09329_ ( .A(fanout_net_21 ), .B(_01322_ ), .C1(_01323_ ), .C2(\u_reg.rf[1][29] ), .ZN(_02198_ ) );
OAI21_X1 _09330_ ( .A(_02198_ ), .B1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01325_ ), .ZN(_02199_ ) );
NAND4_X1 _09331_ ( .A1(_01577_ ), .A2(fanout_net_21 ), .A3(_01322_ ), .A4(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02200_ ) );
NAND3_X1 _09332_ ( .A1(_02199_ ), .A2(_01327_ ), .A3(_02200_ ), .ZN(_02201_ ) );
AND2_X1 _09333_ ( .A1(_02201_ ), .A2(_01046_ ), .ZN(_02202_ ) );
AOI22_X1 _09334_ ( .A1(_01485_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01333_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02203_ ) );
AOI22_X1 _09335_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02204_ ) );
NAND3_X1 _09336_ ( .A1(_02203_ ), .A2(_02204_ ), .A3(_01585_ ), .ZN(_02205_ ) );
AOI21_X1 _09337_ ( .A(_02197_ ), .B1(_02202_ ), .B2(_02205_ ), .ZN(_02206_ ) );
OAI21_X1 _09338_ ( .A(_00736_ ), .B1(_01304_ ), .B2(_02206_ ), .ZN(_02207_ ) );
OR3_X1 _09339_ ( .A1(_02190_ ), .A2(_00723_ ), .A3(_02207_ ), .ZN(_02208_ ) );
NAND4_X1 _09340_ ( .A1(_01416_ ), .A2(_00816_ ), .A3(_00815_ ), .A4(_01538_ ), .ZN(_02209_ ) );
BUF_X4 _09341_ ( .A(_01430_ ), .Z(_02210_ ) );
NAND3_X1 _09342_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][29] ), .A3(_02210_ ), .ZN(_02211_ ) );
NAND3_X1 _09343_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][29] ), .A3(_01435_ ), .ZN(_02212_ ) );
NAND4_X1 _09344_ ( .A1(_01430_ ), .A2(\u_csr.csr[2][29] ), .A3(_01439_ ), .A4(_01442_ ), .ZN(_02213_ ) );
NAND4_X1 _09345_ ( .A1(_01545_ ), .A2(_02211_ ), .A3(_02212_ ), .A4(_02213_ ), .ZN(_02214_ ) );
NAND3_X1 _09346_ ( .A1(_01424_ ), .A2(_01425_ ), .A3(_02214_ ), .ZN(_02215_ ) );
AOI21_X1 _09347_ ( .A(_01535_ ), .B1(_02209_ ), .B2(_02215_ ), .ZN(_02216_ ) );
AOI221_X4 _09348_ ( .A(_02216_ ), .B1(\de_pc[29] ), .B2(_01455_ ), .C1(_01063_ ), .C2(_01065_ ), .ZN(_02217_ ) );
OR3_X1 _09349_ ( .A1(_02190_ ), .A2(_01460_ ), .A3(_02207_ ), .ZN(_02218_ ) );
AOI21_X1 _09350_ ( .A(_01562_ ), .B1(\u_idu.imm_auipc_lui[29] ), .B2(_01563_ ), .ZN(_02219_ ) );
NOR3_X1 _09351_ ( .A1(_02219_ ), .A2(_01555_ ), .A3(_01566_ ), .ZN(_02220_ ) );
AOI211_X1 _09352_ ( .A(_02220_ ), .B(_01053_ ), .C1(\de_pc[29] ), .C2(_01464_ ), .ZN(_02221_ ) );
AOI221_X1 _09353_ ( .A(_01644_ ), .B1(_02208_ ), .B2(_02217_ ), .C1(_02218_ ), .C2(_02221_ ), .ZN(_00141_ ) );
AOI21_X1 _09354_ ( .A(_01884_ ), .B1(_01727_ ), .B2(_01728_ ), .ZN(_02222_ ) );
AOI21_X1 _09355_ ( .A(_01256_ ), .B1(_01732_ ), .B2(_01733_ ), .ZN(_02223_ ) );
MUX2_X1 _09356_ ( .A(\u_lsu.u_clint.mtime[43] ), .B(\u_lsu.u_clint.mtime[11] ), .S(_01209_ ), .Z(_02224_ ) );
AND4_X1 _09357_ ( .A1(\u_lsu.rvalid_clint ), .A2(_01192_ ), .A3(_01211_ ), .A4(_02224_ ), .ZN(_02225_ ) );
AOI21_X1 _09358_ ( .A(_02225_ ), .B1(_01601_ ), .B2(\io_master_rdata[11] ), .ZN(_02226_ ) );
NOR2_X1 _09359_ ( .A1(_02226_ ), .A2(_01253_ ), .ZN(_02227_ ) );
OR3_X1 _09360_ ( .A1(_02222_ ), .A2(_02223_ ), .A3(_02227_ ), .ZN(_02228_ ) );
AOI21_X1 _09361_ ( .A(_01294_ ), .B1(_02059_ ), .B2(_02228_ ), .ZN(_02229_ ) );
NAND2_X1 _09362_ ( .A1(_02229_ ), .A2(fanout_net_12 ), .ZN(_02230_ ) );
MUX2_X1 _09363_ ( .A(\ea_addr[11] ), .B(\u_exu.ecsr[11] ), .S(_01527_ ), .Z(_02231_ ) );
OR2_X1 _09364_ ( .A1(_02231_ ), .A2(fanout_net_12 ), .ZN(_02232_ ) );
AOI21_X1 _09365_ ( .A(_01246_ ), .B1(_02230_ ), .B2(_02232_ ), .ZN(_02233_ ) );
AOI22_X1 _09366_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02234_ ) );
AOI22_X1 _09367_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02235_ ) );
AOI21_X1 _09368_ ( .A(_01318_ ), .B1(_02234_ ), .B2(_02235_ ), .ZN(_02236_ ) );
AOI22_X1 _09369_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02237_ ) );
AOI22_X1 _09370_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02238_ ) );
AOI21_X1 _09371_ ( .A(_01312_ ), .B1(_02237_ ), .B2(_02238_ ), .ZN(_02239_ ) );
OAI21_X1 _09372_ ( .A(_01483_ ), .B1(_02236_ ), .B2(_02239_ ), .ZN(_02240_ ) );
AOI22_X1 _09373_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01495_ ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02241_ ) );
NAND3_X1 _09374_ ( .A1(_01337_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01577_ ), .ZN(_02242_ ) );
NAND3_X1 _09375_ ( .A1(_01337_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01341_ ), .ZN(_02243_ ) );
NAND4_X1 _09376_ ( .A1(_02241_ ), .A2(_01484_ ), .A3(_02242_ ), .A4(_02243_ ), .ZN(_02244_ ) );
NAND3_X1 _09377_ ( .A1(_01337_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01577_ ), .ZN(_02245_ ) );
INV_X1 _09378_ ( .A(\u_reg.rf[1][11] ), .ZN(_02246_ ) );
AOI21_X1 _09379_ ( .A(_01506_ ), .B1(_01341_ ), .B2(_02246_ ), .ZN(_02247_ ) );
NOR2_X1 _09380_ ( .A1(_01341_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02248_ ) );
OAI211_X1 _09381_ ( .A(_01312_ ), .B(_02245_ ), .C1(_02247_ ), .C2(_02248_ ), .ZN(_02249_ ) );
NAND3_X1 _09382_ ( .A1(_02244_ ), .A2(_01046_ ), .A3(_02249_ ), .ZN(_02250_ ) );
AND2_X1 _09383_ ( .A1(_02240_ ), .A2(_02250_ ), .ZN(_02251_ ) );
OAI21_X1 _09384_ ( .A(_00736_ ), .B1(_01304_ ), .B2(_02251_ ), .ZN(_02252_ ) );
OR3_X1 _09385_ ( .A1(_02233_ ), .A2(_00723_ ), .A3(_02252_ ), .ZN(_02253_ ) );
NOR2_X1 _09386_ ( .A1(_01537_ ), .A2(_01419_ ), .ZN(_02254_ ) );
OR2_X1 _09387_ ( .A1(\ea_addr[11] ), .A2(ea_err ), .ZN(_02255_ ) );
OAI211_X1 _09388_ ( .A(_02254_ ), .B(_02255_ ), .C1(_00796_ ), .C2(\ea_pc[11] ), .ZN(_02256_ ) );
AND3_X1 _09389_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][11] ), .A3(_01435_ ), .ZN(_02257_ ) );
AOI21_X1 _09390_ ( .A(_02257_ ), .B1(_01539_ ), .B2(_01783_ ), .ZN(_02258_ ) );
NAND3_X1 _09391_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][11] ), .A3(_02210_ ), .ZN(_02259_ ) );
NAND4_X1 _09392_ ( .A1(_02210_ ), .A2(\u_csr.csr[2][11] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_02260_ ) );
NAND3_X1 _09393_ ( .A1(_02258_ ), .A2(_02259_ ), .A3(_02260_ ), .ZN(_02261_ ) );
NAND3_X1 _09394_ ( .A1(_01776_ ), .A2(_01538_ ), .A3(_02261_ ), .ZN(_02262_ ) );
AOI21_X1 _09395_ ( .A(_01535_ ), .B1(_02256_ ), .B2(_02262_ ), .ZN(_02263_ ) );
AOI221_X4 _09396_ ( .A(_02263_ ), .B1(\de_pc[11] ), .B2(_01455_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_02264_ ) );
OR3_X1 _09397_ ( .A1(_02233_ ), .A2(_01460_ ), .A3(_02252_ ), .ZN(_02265_ ) );
AND3_X1 _09398_ ( .A1(_00665_ ), .A2(\u_idu.imm_branch[11] ), .A3(_00691_ ), .ZN(_02266_ ) );
AOI221_X4 _09399_ ( .A(_02266_ ), .B1(_00726_ ), .B2(\u_idu.imm_auipc_lui[31] ), .C1(fanout_net_22 ), .C2(_00746_ ), .ZN(_02267_ ) );
AND2_X1 _09400_ ( .A1(_01560_ ), .A2(_02267_ ), .ZN(_02268_ ) );
INV_X1 _09401_ ( .A(_02268_ ), .ZN(_02269_ ) );
AOI221_X4 _09402_ ( .A(_01052_ ), .B1(\de_pc[11] ), .B2(_01463_ ), .C1(_01467_ ), .C2(_02269_ ), .ZN(_02270_ ) );
AOI221_X1 _09403_ ( .A(_01644_ ), .B1(_02253_ ), .B2(_02264_ ), .C1(_02265_ ), .C2(_02270_ ), .ZN(_00142_ ) );
AOI22_X1 _09404_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01915_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02271_ ) );
AOI22_X1 _09405_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02272_ ) );
NAND3_X1 _09406_ ( .A1(_02271_ ), .A2(_02272_ ), .A3(_01910_ ), .ZN(_02273_ ) );
AOI22_X1 _09407_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02274_ ) );
AOI22_X1 _09408_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02275_ ) );
NAND3_X1 _09409_ ( .A1(_02274_ ), .A2(_02275_ ), .A3(_01901_ ), .ZN(_02276_ ) );
NAND3_X1 _09410_ ( .A1(_02273_ ), .A2(_02276_ ), .A3(_01756_ ), .ZN(_02277_ ) );
AOI22_X1 _09411_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01915_ ), .B1(_01899_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02278_ ) );
NAND3_X1 _09412_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01903_ ), .ZN(_02279_ ) );
NAND3_X1 _09413_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01905_ ), .ZN(_02280_ ) );
NAND4_X1 _09414_ ( .A1(_02278_ ), .A2(_01901_ ), .A3(_02279_ ), .A4(_02280_ ), .ZN(_02281_ ) );
NAND2_X1 _09415_ ( .A1(_02281_ ), .A2(_01836_ ), .ZN(_02282_ ) );
OAI211_X1 _09416_ ( .A(fanout_net_21 ), .B(_01838_ ), .C1(_01587_ ), .C2(\u_reg.rf[1][10] ), .ZN(_02283_ ) );
OAI21_X1 _09417_ ( .A(_02283_ ), .B1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01905_ ), .ZN(_02284_ ) );
NAND3_X1 _09418_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01903_ ), .ZN(_02285_ ) );
AND3_X1 _09419_ ( .A1(_02284_ ), .A2(_01910_ ), .A3(_02285_ ), .ZN(_02286_ ) );
OAI21_X1 _09420_ ( .A(_02277_ ), .B1(_02282_ ), .B2(_02286_ ), .ZN(_02287_ ) );
AOI21_X1 _09421_ ( .A(_00735_ ), .B1(_01823_ ), .B2(_02287_ ), .ZN(_02288_ ) );
AND3_X1 _09422_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[10] ), .ZN(_02289_ ) );
AOI211_X1 _09423_ ( .A(fanout_net_12 ), .B(_02289_ ), .C1(_01723_ ), .C2(\ea_addr[10] ), .ZN(_02290_ ) );
AND3_X1 _09424_ ( .A1(_01809_ ), .A2(_01270_ ), .A3(_01813_ ), .ZN(_02291_ ) );
AND2_X1 _09425_ ( .A1(_01815_ ), .A2(_01819_ ), .ZN(_02292_ ) );
AOI21_X1 _09426_ ( .A(_02291_ ), .B1(_01255_ ), .B2(_02292_ ), .ZN(_02293_ ) );
NAND2_X1 _09427_ ( .A1(_01598_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ), .ZN(_02294_ ) );
OAI21_X1 _09428_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ), .B1(_01518_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_02295_ ) );
NAND3_X1 _09429_ ( .A1(_02294_ ), .A2(_01670_ ), .A3(_02295_ ), .ZN(_02296_ ) );
NAND3_X1 _09430_ ( .A1(_01192_ ), .A2(_01211_ ), .A3(_02296_ ), .ZN(_02297_ ) );
OAI21_X1 _09431_ ( .A(_02297_ ), .B1(_01681_ ), .B2(\io_master_rdata[10] ), .ZN(_02298_ ) );
OAI21_X1 _09432_ ( .A(_02293_ ), .B1(_01675_ ), .B2(_02298_ ), .ZN(_02299_ ) );
AOI21_X1 _09433_ ( .A(_01295_ ), .B1(_02059_ ), .B2(_02299_ ), .ZN(_02300_ ) );
AOI21_X1 _09434_ ( .A(_02290_ ), .B1(_02300_ ), .B2(fanout_net_12 ), .ZN(\ar_data[10] ) );
OAI21_X1 _09435_ ( .A(_02288_ ), .B1(\ar_data[10] ), .B2(_01825_ ), .ZN(_02301_ ) );
NOR2_X1 _09436_ ( .A1(_02301_ ), .A2(_01770_ ), .ZN(_02302_ ) );
NAND4_X1 _09437_ ( .A1(_01772_ ), .A2(_00814_ ), .A3(_00813_ ), .A4(_01773_ ), .ZN(_02303_ ) );
NAND3_X1 _09438_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][10] ), .A3(_01780_ ), .ZN(_02304_ ) );
AND3_X1 _09439_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][10] ), .A3(_01436_ ), .ZN(_02305_ ) );
AOI21_X1 _09440_ ( .A(_02305_ ), .B1(_01783_ ), .B2(_01626_ ), .ZN(_02306_ ) );
NAND4_X1 _09441_ ( .A1(_01780_ ), .A2(\u_csr.csr[2][10] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_02307_ ) );
NAND3_X1 _09442_ ( .A1(_02304_ ), .A2(_02306_ ), .A3(_02307_ ), .ZN(_02308_ ) );
NAND3_X1 _09443_ ( .A1(_01776_ ), .A2(_01777_ ), .A3(_02308_ ), .ZN(_02309_ ) );
AND2_X1 _09444_ ( .A1(_02303_ ), .A2(_02309_ ), .ZN(_02310_ ) );
INV_X1 _09445_ ( .A(\de_pc[10] ), .ZN(_02311_ ) );
OAI22_X1 _09446_ ( .A1(_02310_ ), .A2(_01791_ ), .B1(_02311_ ), .B2(_01793_ ), .ZN(_02312_ ) );
OAI21_X1 _09447_ ( .A(_01721_ ), .B1(_02302_ ), .B2(_02312_ ), .ZN(_02313_ ) );
OAI22_X1 _09448_ ( .A1(_02301_ ), .A2(_01796_ ), .B1(_02311_ ), .B2(_01797_ ), .ZN(_02314_ ) );
AOI21_X1 _09449_ ( .A(_00862_ ), .B1(_01470_ ), .B2(_00723_ ), .ZN(_02315_ ) );
AND3_X1 _09450_ ( .A1(_00734_ ), .A2(_01121_ ), .A3(_00679_ ), .ZN(_02316_ ) );
NOR2_X1 _09451_ ( .A1(_02315_ ), .A2(_02316_ ), .ZN(_02317_ ) );
INV_X1 _09452_ ( .A(_02317_ ), .ZN(_02318_ ) );
AOI21_X1 _09453_ ( .A(_02314_ ), .B1(_01468_ ), .B2(_02318_ ), .ZN(_02319_ ) );
OAI21_X1 _09454_ ( .A(_02313_ ), .B1(_02319_ ), .B2(_01806_ ), .ZN(_00143_ ) );
AOI21_X1 _09455_ ( .A(_01256_ ), .B1(_01887_ ), .B2(_01888_ ), .ZN(_02320_ ) );
AOI21_X1 _09456_ ( .A(_02320_ ), .B1(_01895_ ), .B2(_01270_ ), .ZN(_02321_ ) );
MUX2_X1 _09457_ ( .A(\u_lsu.u_clint.mtime[41] ), .B(\u_lsu.u_clint.mtime[9] ), .S(_01598_ ), .Z(_02322_ ) );
AND4_X1 _09458_ ( .A1(\u_lsu.rvalid_clint ), .A2(_01666_ ), .A3(_01667_ ), .A4(_02322_ ), .ZN(_02323_ ) );
BUF_X2 _09459_ ( .A(_01601_ ), .Z(io_master_rready ) );
AOI21_X1 _09460_ ( .A(_02323_ ), .B1(io_master_rready ), .B2(\io_master_rdata[9] ), .ZN(_02324_ ) );
OAI21_X1 _09461_ ( .A(_02321_ ), .B1(_01664_ ), .B2(_02324_ ), .ZN(_02325_ ) );
AOI21_X1 _09462_ ( .A(_01294_ ), .B1(_02059_ ), .B2(_02325_ ), .ZN(_02326_ ) );
NAND2_X1 _09463_ ( .A1(_02326_ ), .A2(fanout_net_12 ), .ZN(_02327_ ) );
MUX2_X1 _09464_ ( .A(\ea_addr[9] ), .B(\u_exu.ecsr[9] ), .S(_01298_ ), .Z(_02328_ ) );
OR2_X1 _09465_ ( .A1(_02328_ ), .A2(fanout_net_12 ), .ZN(_02329_ ) );
AOI21_X1 _09466_ ( .A(_01246_ ), .B1(_02327_ ), .B2(_02329_ ), .ZN(_02330_ ) );
AOI22_X1 _09467_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02331_ ) );
AOI22_X1 _09468_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02332_ ) );
NAND3_X1 _09469_ ( .A1(_02331_ ), .A2(_02332_ ), .A3(_01312_ ), .ZN(_02333_ ) );
AOI22_X1 _09470_ ( .A1(_01005_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02334_ ) );
AOI22_X1 _09471_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02335_ ) );
NAND3_X1 _09472_ ( .A1(_02334_ ), .A2(_02335_ ), .A3(_01318_ ), .ZN(_02336_ ) );
AND3_X1 _09473_ ( .A1(_02333_ ), .A2(_02336_ ), .A3(_01320_ ), .ZN(_02337_ ) );
OAI211_X1 _09474_ ( .A(fanout_net_21 ), .B(_01322_ ), .C1(_01323_ ), .C2(\u_reg.rf[1][9] ), .ZN(_02338_ ) );
OAI21_X1 _09475_ ( .A(_02338_ ), .B1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01325_ ), .ZN(_02339_ ) );
NAND4_X1 _09476_ ( .A1(_01577_ ), .A2(fanout_net_21 ), .A3(_01322_ ), .A4(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02340_ ) );
NAND3_X1 _09477_ ( .A1(_02339_ ), .A2(_01327_ ), .A3(_02340_ ), .ZN(_02341_ ) );
AND2_X1 _09478_ ( .A1(_02341_ ), .A2(_01046_ ), .ZN(_02342_ ) );
AOI22_X1 _09479_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01333_ ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02343_ ) );
NAND3_X1 _09480_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01339_ ), .ZN(_02344_ ) );
NAND3_X1 _09481_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01342_ ), .ZN(_02345_ ) );
NAND4_X1 _09482_ ( .A1(_02343_ ), .A2(_01336_ ), .A3(_02344_ ), .A4(_02345_ ), .ZN(_02346_ ) );
AOI21_X1 _09483_ ( .A(_02337_ ), .B1(_02342_ ), .B2(_02346_ ), .ZN(_02347_ ) );
OAI21_X1 _09484_ ( .A(_00736_ ), .B1(_01304_ ), .B2(_02347_ ), .ZN(_02348_ ) );
OR3_X1 _09485_ ( .A1(_02330_ ), .A2(_00723_ ), .A3(_02348_ ), .ZN(_02349_ ) );
NAND4_X1 _09486_ ( .A1(_01416_ ), .A2(_00818_ ), .A3(_00817_ ), .A4(_01421_ ), .ZN(_02350_ ) );
NAND3_X1 _09487_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][9] ), .A3(_01431_ ), .ZN(_02351_ ) );
NAND3_X1 _09488_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][9] ), .A3(_01436_ ), .ZN(_02352_ ) );
NAND4_X1 _09489_ ( .A1(_02210_ ), .A2(\u_csr.csr[2][9] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_02353_ ) );
NAND3_X1 _09490_ ( .A1(_02351_ ), .A2(_02352_ ), .A3(_02353_ ), .ZN(_02354_ ) );
NAND3_X1 _09491_ ( .A1(_01537_ ), .A2(_01538_ ), .A3(_02354_ ), .ZN(_02355_ ) );
AOI21_X1 _09492_ ( .A(_01535_ ), .B1(_02350_ ), .B2(_02355_ ), .ZN(_02356_ ) );
AOI221_X4 _09493_ ( .A(_02356_ ), .B1(\de_pc[9] ), .B2(_01455_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_02357_ ) );
OR3_X1 _09494_ ( .A1(_02330_ ), .A2(_01460_ ), .A3(_02348_ ), .ZN(_02358_ ) );
AOI21_X1 _09495_ ( .A(_00743_ ), .B1(_00679_ ), .B2(_00734_ ), .ZN(_02359_ ) );
AND2_X1 _09496_ ( .A1(_01470_ ), .A2(_02359_ ), .ZN(_02360_ ) );
NOR2_X1 _09497_ ( .A1(_02360_ ), .A2(_00889_ ), .ZN(_02361_ ) );
AOI221_X4 _09498_ ( .A(_01052_ ), .B1(\de_pc[9] ), .B2(_01463_ ), .C1(_01467_ ), .C2(_02361_ ), .ZN(_02362_ ) );
AOI221_X1 _09499_ ( .A(_01644_ ), .B1(_02349_ ), .B2(_02357_ ), .C1(_02358_ ), .C2(_02362_ ), .ZN(_00144_ ) );
AND3_X1 _09500_ ( .A1(\ea_mask[0] ), .A2(\u_exu.eopt[15] ), .A3(\u_exu.ecsr[8] ), .ZN(_02363_ ) );
AOI211_X1 _09501_ ( .A(fanout_net_12 ), .B(_02363_ ), .C1(_01723_ ), .C2(\ea_addr[8] ), .ZN(_02364_ ) );
NAND3_X1 _09502_ ( .A1(_01945_ ), .A2(_01270_ ), .A3(_01951_ ), .ZN(_02365_ ) );
OAI211_X1 _09503_ ( .A(_01255_ ), .B(_01958_ ), .C1(_01681_ ), .C2(\io_master_rdata[24] ), .ZN(_02366_ ) );
AND2_X1 _09504_ ( .A1(_02365_ ), .A2(_02366_ ), .ZN(_02367_ ) );
INV_X1 _09505_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ), .ZN(_02368_ ) );
OR3_X1 _09506_ ( .A1(_01946_ ), .A2(\u_arbiter.raddr[2] ), .A3(_02368_ ), .ZN(_02369_ ) );
OAI21_X1 _09507_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ), .B1(_01946_ ), .B2(\u_arbiter.raddr[2] ), .ZN(_02370_ ) );
NAND3_X1 _09508_ ( .A1(_02369_ ), .A2(_01670_ ), .A3(_02370_ ), .ZN(_02371_ ) );
NAND3_X1 _09509_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(_02371_ ), .ZN(_02372_ ) );
OAI21_X1 _09510_ ( .A(_02372_ ), .B1(_01681_ ), .B2(\io_master_rdata[8] ), .ZN(_02373_ ) );
OAI21_X1 _09511_ ( .A(_02367_ ), .B1(_01675_ ), .B2(_02373_ ), .ZN(_02374_ ) );
AOI21_X1 _09512_ ( .A(_01295_ ), .B1(_02059_ ), .B2(_02374_ ), .ZN(_02375_ ) );
AOI21_X2 _09513_ ( .A(_02364_ ), .B1(_02375_ ), .B2(fanout_net_12 ), .ZN(\ar_data[8] ) );
NOR2_X1 _09514_ ( .A1(\ar_data[8] ), .A2(_01246_ ), .ZN(_02376_ ) );
AOI22_X1 _09515_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02377_ ) );
AOI22_X1 _09516_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02378_ ) );
NAND3_X1 _09517_ ( .A1(_02377_ ), .A2(_02378_ ), .A3(_01585_ ), .ZN(_02379_ ) );
OAI211_X1 _09518_ ( .A(fanout_net_21 ), .B(_01837_ ), .C1(_01339_ ), .C2(\u_reg.rf[1][8] ), .ZN(_02380_ ) );
OAI21_X1 _09519_ ( .A(_02380_ ), .B1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01750_ ), .ZN(_02381_ ) );
NAND4_X1 _09520_ ( .A1(_01587_ ), .A2(fanout_net_21 ), .A3(_01837_ ), .A4(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02382_ ) );
NAND3_X1 _09521_ ( .A1(_02381_ ), .A2(_01746_ ), .A3(_02382_ ), .ZN(_02383_ ) );
NAND3_X1 _09522_ ( .A1(_02379_ ), .A2(_01504_ ), .A3(_02383_ ), .ZN(_02384_ ) );
AOI22_X1 _09523_ ( .A1(_01485_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01333_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02385_ ) );
AOI22_X1 _09524_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02386_ ) );
AOI21_X1 _09525_ ( .A(_01585_ ), .B1(_02385_ ), .B2(_02386_ ), .ZN(_02387_ ) );
AOI22_X1 _09526_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02388_ ) );
AOI22_X1 _09527_ ( .A1(_01485_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01486_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02389_ ) );
AOI21_X1 _09528_ ( .A(_01580_ ), .B1(_02388_ ), .B2(_02389_ ), .ZN(_02390_ ) );
OAI21_X1 _09529_ ( .A(_01483_ ), .B1(_02387_ ), .B2(_02390_ ), .ZN(_02391_ ) );
AOI21_X1 _09530_ ( .A(_01244_ ), .B1(_02384_ ), .B2(_02391_ ), .ZN(_02392_ ) );
NOR3_X4 _09531_ ( .A1(_02376_ ), .A2(_00735_ ), .A3(_02392_ ), .ZN(_02393_ ) );
NAND2_X1 _09532_ ( .A1(_02393_ ), .A2(_01533_ ), .ZN(_02394_ ) );
NAND4_X1 _09533_ ( .A1(_01416_ ), .A2(_00820_ ), .A3(_00819_ ), .A4(_01538_ ), .ZN(_02395_ ) );
AND3_X1 _09534_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][8] ), .A3(_01435_ ), .ZN(_02396_ ) );
AOI21_X1 _09535_ ( .A(_02396_ ), .B1(_01928_ ), .B2(_01783_ ), .ZN(_02397_ ) );
NAND3_X1 _09536_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][8] ), .A3(_01431_ ), .ZN(_02398_ ) );
NAND4_X1 _09537_ ( .A1(_01431_ ), .A2(\u_csr.csr[2][8] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_02399_ ) );
NAND3_X1 _09538_ ( .A1(_02397_ ), .A2(_02398_ ), .A3(_02399_ ), .ZN(_02400_ ) );
NAND3_X1 _09539_ ( .A1(_01776_ ), .A2(_01425_ ), .A3(_02400_ ), .ZN(_02401_ ) );
AOI21_X1 _09540_ ( .A(_01535_ ), .B1(_02395_ ), .B2(_02401_ ), .ZN(_02402_ ) );
AOI221_X4 _09541_ ( .A(_02402_ ), .B1(\de_pc[8] ), .B2(_01454_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_02403_ ) );
NAND2_X1 _09542_ ( .A1(_02393_ ), .A2(_01556_ ), .ZN(_02404_ ) );
NOR2_X1 _09543_ ( .A1(_02360_ ), .A2(_00890_ ), .ZN(_02405_ ) );
AOI221_X4 _09544_ ( .A(_01052_ ), .B1(\de_pc[8] ), .B2(_01463_ ), .C1(_01467_ ), .C2(_02405_ ), .ZN(_02406_ ) );
AOI221_X1 _09545_ ( .A(_01644_ ), .B1(_02394_ ), .B2(_02403_ ), .C1(_02404_ ), .C2(_02406_ ), .ZN(_00145_ ) );
BUF_X4 _09546_ ( .A(_01466_ ), .Z(_02407_ ) );
NOR2_X1 _09547_ ( .A1(_02360_ ), .A2(_00707_ ), .ZN(_02408_ ) );
NAND3_X1 _09548_ ( .A1(_01460_ ), .A2(_02407_ ), .A3(_02408_ ), .ZN(_02409_ ) );
INV_X1 _09549_ ( .A(\de_pc[7] ), .ZN(_02410_ ) );
MUX2_X1 _09550_ ( .A(\ea_addr[7] ), .B(\u_exu.ecsr[7] ), .S(_01299_ ), .Z(_02411_ ) );
AND2_X2 _09551_ ( .A1(_01273_ ), .A2(_01292_ ), .ZN(_02412_ ) );
NOR2_X1 _09552_ ( .A1(_01291_ ), .A2(_02412_ ), .ZN(_02413_ ) );
MUX2_X1 _09553_ ( .A(_02411_ ), .B(_02413_ ), .S(fanout_net_12 ), .Z(\ar_data[7] ) );
NOR2_X1 _09554_ ( .A1(\ar_data[7] ), .A2(_01823_ ), .ZN(_02414_ ) );
AOI22_X1 _09555_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01915_ ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02415_ ) );
NAND3_X1 _09556_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01903_ ), .ZN(_02416_ ) );
NAND3_X1 _09557_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01905_ ), .ZN(_02417_ ) );
NAND4_X1 _09558_ ( .A1(_02415_ ), .A2(_01744_ ), .A3(_02416_ ), .A4(_02417_ ), .ZN(_02418_ ) );
NAND3_X1 _09559_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01748_ ), .ZN(_02419_ ) );
INV_X1 _09560_ ( .A(\u_reg.rf[1][7] ), .ZN(_02420_ ) );
AOI21_X1 _09561_ ( .A(_01506_ ), .B1(_01905_ ), .B2(_02420_ ), .ZN(_02421_ ) );
NOR2_X1 _09562_ ( .A1(_01905_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02422_ ) );
OAI211_X1 _09563_ ( .A(_01746_ ), .B(_02419_ ), .C1(_02421_ ), .C2(_02422_ ), .ZN(_02423_ ) );
NAND3_X1 _09564_ ( .A1(_02418_ ), .A2(_01836_ ), .A3(_02423_ ), .ZN(_02424_ ) );
AOI22_X1 _09565_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02425_ ) );
AOI22_X1 _09566_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02426_ ) );
NAND3_X1 _09567_ ( .A1(_02425_ ), .A2(_02426_ ), .A3(_01910_ ), .ZN(_02427_ ) );
AOI22_X1 _09568_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01742_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02428_ ) );
AOI22_X1 _09569_ ( .A1(_01738_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01739_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02429_ ) );
NAND3_X1 _09570_ ( .A1(_02428_ ), .A2(_02429_ ), .A3(_01744_ ), .ZN(_02430_ ) );
NAND3_X1 _09571_ ( .A1(_02427_ ), .A2(_02430_ ), .A3(_01756_ ), .ZN(_02431_ ) );
AOI21_X1 _09572_ ( .A(_01482_ ), .B1(_02424_ ), .B2(_02431_ ), .ZN(_02432_ ) );
OR3_X1 _09573_ ( .A1(_02414_ ), .A2(_01999_ ), .A3(_02432_ ), .ZN(_02433_ ) );
OAI221_X1 _09574_ ( .A(_02409_ ), .B1(_02410_ ), .B2(_01797_ ), .C1(_02433_ ), .C2(_01796_ ), .ZN(_02434_ ) );
NAND2_X1 _09575_ ( .A1(_02434_ ), .A2(_01078_ ), .ZN(_02435_ ) );
NOR2_X1 _09576_ ( .A1(_02433_ ), .A2(_01770_ ), .ZN(_02436_ ) );
AND4_X1 _09577_ ( .A1(_00822_ ), .A2(_01772_ ), .A3(_00821_ ), .A4(_01777_ ), .ZN(_02437_ ) );
NAND3_X1 _09578_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][7] ), .A3(_01779_ ), .ZN(_02438_ ) );
NAND3_X1 _09579_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][7] ), .A3(_01874_ ), .ZN(_02439_ ) );
NAND4_X1 _09580_ ( .A1(_01779_ ), .A2(\u_csr.csr[2][7] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_02440_ ) );
NAND4_X1 _09581_ ( .A1(_01692_ ), .A2(_02438_ ), .A3(_02439_ ), .A4(_02440_ ), .ZN(_02441_ ) );
AND3_X1 _09582_ ( .A1(_01424_ ), .A2(_01777_ ), .A3(_02441_ ), .ZN(_02442_ ) );
OAI21_X1 _09583_ ( .A(_01351_ ), .B1(_02437_ ), .B2(_02442_ ), .ZN(_02443_ ) );
OAI21_X1 _09584_ ( .A(_02443_ ), .B1(_02410_ ), .B2(_01793_ ), .ZN(_02444_ ) );
OAI21_X1 _09585_ ( .A(_01053_ ), .B1(_02436_ ), .B2(_02444_ ), .ZN(_02445_ ) );
AOI21_X1 _09586_ ( .A(_01076_ ), .B1(_02435_ ), .B2(_02445_ ), .ZN(_00146_ ) );
AOI22_X1 _09587_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02446_ ) );
AOI22_X1 _09588_ ( .A1(_01741_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02447_ ) );
NAND3_X1 _09589_ ( .A1(_02446_ ), .A2(_02447_ ), .A3(_01746_ ), .ZN(_02448_ ) );
AOI22_X1 _09590_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02449_ ) );
AOI22_X1 _09591_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02450_ ) );
NAND3_X1 _09592_ ( .A1(_02449_ ), .A2(_02450_ ), .A3(_01744_ ), .ZN(_02451_ ) );
NAND3_X1 _09593_ ( .A1(_02448_ ), .A2(_02451_ ), .A3(_01756_ ), .ZN(_02452_ ) );
OAI211_X1 _09594_ ( .A(fanout_net_21 ), .B(_01837_ ), .C1(_01587_ ), .C2(\u_reg.rf[1][6] ), .ZN(_02453_ ) );
OAI21_X1 _09595_ ( .A(_02453_ ), .B1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01750_ ), .ZN(_02454_ ) );
NAND3_X1 _09596_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01748_ ), .ZN(_02455_ ) );
AND3_X1 _09597_ ( .A1(_02454_ ), .A2(_01746_ ), .A3(_02455_ ), .ZN(_02456_ ) );
AOI22_X1 _09598_ ( .A1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01739_ ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02457_ ) );
NAND3_X1 _09599_ ( .A1(_01747_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01748_ ), .ZN(_02458_ ) );
NAND3_X1 _09600_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01750_ ), .ZN(_02459_ ) );
NAND4_X1 _09601_ ( .A1(_02457_ ), .A2(_01744_ ), .A3(_02458_ ), .A4(_02459_ ), .ZN(_02460_ ) );
NAND2_X1 _09602_ ( .A1(_02460_ ), .A2(_01504_ ), .ZN(_02461_ ) );
OAI211_X1 _09603_ ( .A(_01246_ ), .B(_02452_ ), .C1(_02456_ ), .C2(_02461_ ), .ZN(_02462_ ) );
MUX2_X1 _09604_ ( .A(\ea_addr[6] ), .B(\u_exu.ecsr[6] ), .S(_01527_ ), .Z(_02463_ ) );
NOR2_X1 _09605_ ( .A1(_02463_ ), .A2(fanout_net_12 ), .ZN(_02464_ ) );
INV_X1 _09606_ ( .A(_02412_ ), .ZN(_02465_ ) );
INV_X1 _09607_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ), .ZN(_02466_ ) );
OR3_X1 _09608_ ( .A1(_01946_ ), .A2(\u_arbiter.raddr[2] ), .A3(_02466_ ), .ZN(_02467_ ) );
NAND2_X1 _09609_ ( .A1(_02467_ ), .A2(_01670_ ), .ZN(_02468_ ) );
AOI211_X1 _09610_ ( .A(_02468_ ), .B(io_master_rready ), .C1(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ), .C2(_02116_ ), .ZN(_02469_ ) );
AOI21_X1 _09611_ ( .A(_02469_ ), .B1(io_master_rready ), .B2(\io_master_rdata[6] ), .ZN(_02470_ ) );
NOR2_X1 _09612_ ( .A1(_02470_ ), .A2(_01675_ ), .ZN(_02471_ ) );
AND3_X1 _09613_ ( .A1(_01514_ ), .A2(_01281_ ), .A3(_01521_ ), .ZN(_02472_ ) );
AOI21_X1 _09614_ ( .A(_02472_ ), .B1(_01255_ ), .B2(_02067_ ), .ZN(_02473_ ) );
OAI21_X1 _09615_ ( .A(_02473_ ), .B1(_01884_ ), .B2(_02073_ ), .ZN(_02474_ ) );
OAI21_X1 _09616_ ( .A(_02465_ ), .B1(_02471_ ), .B2(_02474_ ), .ZN(_02475_ ) );
AOI21_X1 _09617_ ( .A(_02464_ ), .B1(_02475_ ), .B2(fanout_net_12 ), .ZN(\ar_data[6] ) );
NAND3_X1 _09618_ ( .A1(\ar_data[6] ), .A2(_01223_ ), .A3(_01243_ ), .ZN(_02476_ ) );
AOI21_X1 _09619_ ( .A(_00735_ ), .B1(_02462_ ), .B2(_02476_ ), .ZN(_02477_ ) );
NAND2_X1 _09620_ ( .A1(_02477_ ), .A2(_01533_ ), .ZN(_02478_ ) );
AND4_X1 _09621_ ( .A1(\u_csr.csr[2][6] ), .A2(_01539_ ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_02479_ ) );
NOR3_X1 _09622_ ( .A1(_02479_ ), .A2(_01544_ ), .A3(_01627_ ), .ZN(_02480_ ) );
AND4_X1 _09623_ ( .A1(\u_csr.csr[0][6] ), .A2(_01439_ ), .A3(_01410_ ), .A4(_01548_ ), .ZN(_02481_ ) );
AOI21_X1 _09624_ ( .A(_02481_ ), .B1(_01631_ ), .B2(\u_csr.csr[1][6] ), .ZN(_02482_ ) );
AOI21_X1 _09625_ ( .A(_01619_ ), .B1(_02480_ ), .B2(_02482_ ), .ZN(_02483_ ) );
AOI211_X1 _09626_ ( .A(_01419_ ), .B(_01537_ ), .C1(_00823_ ), .C2(_00824_ ), .ZN(_02484_ ) );
NOR2_X1 _09627_ ( .A1(_02483_ ), .A2(_02484_ ), .ZN(_02485_ ) );
NOR2_X1 _09628_ ( .A1(_02485_ ), .A2(_01353_ ), .ZN(_02486_ ) );
AOI211_X1 _09629_ ( .A(_01077_ ), .B(_02486_ ), .C1(\de_pc[6] ), .C2(_01455_ ), .ZN(_02487_ ) );
NAND2_X1 _09630_ ( .A1(_02477_ ), .A2(_01556_ ), .ZN(_02488_ ) );
NOR2_X1 _09631_ ( .A1(_02360_ ), .A2(_00880_ ), .ZN(_02489_ ) );
AOI221_X4 _09632_ ( .A(_01051_ ), .B1(\de_pc[6] ), .B2(_01463_ ), .C1(_01467_ ), .C2(_02489_ ), .ZN(_02490_ ) );
AOI221_X4 _09633_ ( .A(_01644_ ), .B1(_02478_ ), .B2(_02487_ ), .C1(_02488_ ), .C2(_02490_ ), .ZN(_00147_ ) );
MUX2_X1 _09634_ ( .A(\ea_addr[5] ), .B(\u_exu.ecsr[5] ), .S(_01299_ ), .Z(_02491_ ) );
OR2_X1 _09635_ ( .A1(_01608_ ), .A2(_01282_ ), .ZN(_02492_ ) );
NOR2_X1 _09636_ ( .A1(_02118_ ), .A2(_01884_ ), .ZN(_02493_ ) );
AOI21_X1 _09637_ ( .A(_01256_ ), .B1(_01600_ ), .B2(_01602_ ), .ZN(_02494_ ) );
NOR2_X1 _09638_ ( .A1(_02493_ ), .A2(_02494_ ), .ZN(_02495_ ) );
AND3_X1 _09639_ ( .A1(_02492_ ), .A2(_01664_ ), .A3(_02495_ ), .ZN(_02496_ ) );
OR3_X1 _09640_ ( .A1(_01946_ ), .A2(\u_arbiter.raddr[2] ), .A3(\u_lsu.u_clint.mtime[5] ), .ZN(_02497_ ) );
OAI211_X1 _09641_ ( .A(_01595_ ), .B(_02497_ ), .C1(\u_lsu.u_clint.mtime[37] ), .C2(_01599_ ), .ZN(_02498_ ) );
AOI21_X1 _09642_ ( .A(_01664_ ), .B1(io_master_rready ), .B2(\io_master_rdata[5] ), .ZN(_02499_ ) );
AND2_X1 _09643_ ( .A1(_02498_ ), .A2(_02499_ ), .ZN(_02500_ ) );
NOR3_X1 _09644_ ( .A1(_02496_ ), .A2(_02412_ ), .A3(_02500_ ), .ZN(_02501_ ) );
MUX2_X1 _09645_ ( .A(_02491_ ), .B(_02501_ ), .S(fanout_net_12 ), .Z(\ar_data[5] ) );
NAND2_X1 _09646_ ( .A1(\ar_data[5] ), .A2(_01482_ ), .ZN(_02502_ ) );
AOI22_X1 _09647_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02503_ ) );
AOI22_X1 _09648_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02504_ ) );
NAND3_X1 _09649_ ( .A1(_02503_ ), .A2(_02504_ ), .A3(_01746_ ), .ZN(_02505_ ) );
AOI22_X1 _09650_ ( .A1(_01760_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01761_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02506_ ) );
AOI22_X1 _09651_ ( .A1(_01757_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02507_ ) );
NAND3_X1 _09652_ ( .A1(_02506_ ), .A2(_02507_ ), .A3(_01585_ ), .ZN(_02508_ ) );
NAND3_X1 _09653_ ( .A1(_02505_ ), .A2(_02508_ ), .A3(_01756_ ), .ZN(_02509_ ) );
AOI22_X1 _09654_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01758_ ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02510_ ) );
NAND3_X1 _09655_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01748_ ), .ZN(_02511_ ) );
NAND3_X1 _09656_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01750_ ), .ZN(_02512_ ) );
AND4_X1 _09657_ ( .A1(_01744_ ), .A2(_02510_ ), .A3(_02511_ ), .A4(_02512_ ), .ZN(_02513_ ) );
OAI21_X1 _09658_ ( .A(_00976_ ), .B1(_01341_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02514_ ) );
OAI21_X1 _09659_ ( .A(_02514_ ), .B1(\u_reg.rf[1][5] ), .B2(_01328_ ), .ZN(_02515_ ) );
AOI211_X1 _09660_ ( .A(_01336_ ), .B(_02515_ ), .C1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_01757_ ), .ZN(_02516_ ) );
OR2_X1 _09661_ ( .A1(_02516_ ), .A2(_01483_ ), .ZN(_02517_ ) );
OAI211_X1 _09662_ ( .A(_01246_ ), .B(_02509_ ), .C1(_02513_ ), .C2(_02517_ ), .ZN(_02518_ ) );
AOI21_X1 _09663_ ( .A(_00735_ ), .B1(_02502_ ), .B2(_02518_ ), .ZN(_02519_ ) );
NAND2_X1 _09664_ ( .A1(_02519_ ), .A2(_00743_ ), .ZN(_02520_ ) );
AND4_X1 _09665_ ( .A1(\u_csr.csr[2][5] ), .A2(_01539_ ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_02521_ ) );
NOR3_X1 _09666_ ( .A1(_02521_ ), .A2(_01544_ ), .A3(_01627_ ), .ZN(_02522_ ) );
AND4_X1 _09667_ ( .A1(\u_csr.csr[0][5] ), .A2(_01439_ ), .A3(_01410_ ), .A4(_01548_ ), .ZN(_02523_ ) );
AOI21_X1 _09668_ ( .A(_02523_ ), .B1(_01631_ ), .B2(\u_csr.csr[1][5] ), .ZN(_02524_ ) );
AOI21_X1 _09669_ ( .A(_01619_ ), .B1(_02522_ ), .B2(_02524_ ), .ZN(_02525_ ) );
AOI211_X1 _09670_ ( .A(_01419_ ), .B(_01537_ ), .C1(_00825_ ), .C2(_00826_ ), .ZN(_02526_ ) );
NOR2_X1 _09671_ ( .A1(_02525_ ), .A2(_02526_ ), .ZN(_02527_ ) );
NOR2_X1 _09672_ ( .A1(_02527_ ), .A2(_01353_ ), .ZN(_02528_ ) );
AOI211_X1 _09673_ ( .A(_01077_ ), .B(_02528_ ), .C1(\de_pc[5] ), .C2(_01455_ ), .ZN(_02529_ ) );
NAND2_X1 _09674_ ( .A1(_02519_ ), .A2(_01556_ ), .ZN(_02530_ ) );
NOR2_X1 _09675_ ( .A1(_02360_ ), .A2(_00891_ ), .ZN(_02531_ ) );
AOI221_X4 _09676_ ( .A(_01051_ ), .B1(\de_pc[5] ), .B2(_01463_ ), .C1(_01467_ ), .C2(_02531_ ), .ZN(_02532_ ) );
AOI221_X4 _09677_ ( .A(_01644_ ), .B1(_02520_ ), .B2(_02529_ ), .C1(_02530_ ), .C2(_02532_ ), .ZN(_00148_ ) );
AOI22_X1 _09678_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01826_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02533_ ) );
AOI22_X1 _09679_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02534_ ) );
NAND3_X1 _09680_ ( .A1(_02533_ ), .A2(_02534_ ), .A3(_01841_ ), .ZN(_02535_ ) );
AOI22_X1 _09681_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02536_ ) );
AOI22_X1 _09682_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02537_ ) );
NAND3_X1 _09683_ ( .A1(_02536_ ), .A2(_02537_ ), .A3(_01829_ ), .ZN(_02538_ ) );
NAND3_X1 _09684_ ( .A1(_02535_ ), .A2(_02538_ ), .A3(_01855_ ), .ZN(_02539_ ) );
OAI211_X1 _09685_ ( .A(fanout_net_21 ), .B(_01838_ ), .C1(_01903_ ), .C2(\u_reg.rf[1][4] ), .ZN(_02540_ ) );
OAI21_X1 _09686_ ( .A(_02540_ ), .B1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01833_ ), .ZN(_02541_ ) );
NAND3_X1 _09687_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_02542_ ) );
AND3_X1 _09688_ ( .A1(_02541_ ), .A2(_01841_ ), .A3(_02542_ ), .ZN(_02543_ ) );
AOI22_X1 _09689_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01826_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02544_ ) );
AOI22_X1 _09690_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02545_ ) );
NAND3_X1 _09691_ ( .A1(_02544_ ), .A2(_02545_ ), .A3(_01829_ ), .ZN(_02546_ ) );
NAND2_X1 _09692_ ( .A1(_02546_ ), .A2(_01836_ ), .ZN(_02547_ ) );
OAI211_X1 _09693_ ( .A(_01823_ ), .B(_02539_ ), .C1(_02543_ ), .C2(_02547_ ), .ZN(_02548_ ) );
NOR2_X1 _09694_ ( .A1(_02166_ ), .A2(_01884_ ), .ZN(_02549_ ) );
INV_X1 _09695_ ( .A(_02549_ ), .ZN(_02550_ ) );
AND3_X1 _09696_ ( .A1(_01665_ ), .A2(_01255_ ), .A3(_01673_ ), .ZN(_02551_ ) );
AOI21_X1 _09697_ ( .A(_02551_ ), .B1(_01281_ ), .B2(_02160_ ), .ZN(_02552_ ) );
AND3_X1 _09698_ ( .A1(_02550_ ), .A2(_02552_ ), .A3(_01664_ ), .ZN(_02553_ ) );
INV_X1 _09699_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_26_A_$_ANDNOT__Y_B ), .ZN(_02554_ ) );
NOR2_X1 _09700_ ( .A1(_01599_ ), .A2(_02554_ ), .ZN(_02555_ ) );
AND2_X1 _09701_ ( .A1(_01598_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ), .ZN(_02556_ ) );
NOR4_X1 _09702_ ( .A1(_01601_ ), .A2(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .A3(_02555_ ), .A4(_02556_ ), .ZN(_02557_ ) );
AOI21_X1 _09703_ ( .A(_02557_ ), .B1(io_master_rready ), .B2(\io_master_rdata[4] ), .ZN(_02558_ ) );
AND2_X1 _09704_ ( .A1(_02558_ ), .A2(_01523_ ), .ZN(_02559_ ) );
NOR3_X1 _09705_ ( .A1(_02553_ ), .A2(_02412_ ), .A3(_02559_ ), .ZN(_02560_ ) );
OR2_X1 _09706_ ( .A1(_02560_ ), .A2(_01129_ ), .ZN(_02561_ ) );
MUX2_X1 _09707_ ( .A(\ea_addr[4] ), .B(\u_exu.ecsr[4] ), .S(_01299_ ), .Z(_02562_ ) );
OR2_X1 _09708_ ( .A1(_02562_ ), .A2(fanout_net_12 ), .ZN(_02563_ ) );
NAND3_X1 _09709_ ( .A1(_02561_ ), .A2(_01531_ ), .A3(_02563_ ), .ZN(_02564_ ) );
AOI21_X1 _09710_ ( .A(_01999_ ), .B1(_02548_ ), .B2(_02564_ ), .ZN(_02565_ ) );
AND2_X1 _09711_ ( .A1(_02565_ ), .A2(_01533_ ), .ZN(_02566_ ) );
NAND4_X1 _09712_ ( .A1(_01772_ ), .A2(_00828_ ), .A3(_00827_ ), .A4(_01425_ ), .ZN(_02567_ ) );
NAND3_X1 _09713_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][4] ), .A3(_01779_ ), .ZN(_02568_ ) );
NAND3_X1 _09714_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][4] ), .A3(_01874_ ), .ZN(_02569_ ) );
NAND4_X1 _09715_ ( .A1(_01779_ ), .A2(\u_csr.csr[2][4] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_02570_ ) );
NAND4_X1 _09716_ ( .A1(_01545_ ), .A2(_02568_ ), .A3(_02569_ ), .A4(_02570_ ), .ZN(_02571_ ) );
NAND3_X1 _09717_ ( .A1(_01424_ ), .A2(_01773_ ), .A3(_02571_ ), .ZN(_02572_ ) );
AND2_X1 _09718_ ( .A1(_02567_ ), .A2(_02572_ ), .ZN(_02573_ ) );
INV_X1 _09719_ ( .A(\de_pc[4] ), .ZN(_02574_ ) );
OAI22_X1 _09720_ ( .A1(_02573_ ), .A2(_01791_ ), .B1(_02574_ ), .B2(_01453_ ), .ZN(_02575_ ) );
OAI21_X1 _09721_ ( .A(_01721_ ), .B1(_02566_ ), .B2(_02575_ ), .ZN(_02576_ ) );
NAND2_X1 _09722_ ( .A1(_02565_ ), .A2(_01557_ ), .ZN(_02577_ ) );
BUF_X4 _09723_ ( .A(_01460_ ), .Z(_02578_ ) );
AOI21_X1 _09724_ ( .A(_00734_ ), .B1(_00687_ ), .B2(_00720_ ), .ZN(_02579_ ) );
AND2_X1 _09725_ ( .A1(_02579_ ), .A2(_00924_ ), .ZN(_02580_ ) );
OR2_X1 _09726_ ( .A1(_02580_ ), .A2(_00892_ ), .ZN(_02581_ ) );
OAI21_X1 _09727_ ( .A(\u_idu.imm_branch[4] ), .B1(_00727_ ), .B2(_00692_ ), .ZN(_02582_ ) );
NAND2_X1 _09728_ ( .A1(_02581_ ), .A2(_02582_ ), .ZN(_02583_ ) );
NAND3_X1 _09729_ ( .A1(_02578_ ), .A2(_02407_ ), .A3(_02583_ ), .ZN(_02584_ ) );
NAND3_X1 _09730_ ( .A1(_02578_ ), .A2(\de_pc[4] ), .A3(_01861_ ), .ZN(_02585_ ) );
AND3_X1 _09731_ ( .A1(_02577_ ), .A2(_02584_ ), .A3(_02585_ ), .ZN(_02586_ ) );
OAI21_X1 _09732_ ( .A(_02576_ ), .B1(_02586_ ), .B2(_01806_ ), .ZN(_00149_ ) );
MUX2_X1 _09733_ ( .A(\ea_addr[3] ), .B(\u_exu.ecsr[3] ), .S(_01299_ ), .Z(_02587_ ) );
OR2_X1 _09734_ ( .A1(_01734_ ), .A2(_01282_ ), .ZN(_02588_ ) );
AOI21_X1 _09735_ ( .A(_01256_ ), .B1(_01727_ ), .B2(_01728_ ), .ZN(_02589_ ) );
NOR2_X1 _09736_ ( .A1(_02226_ ), .A2(_01884_ ), .ZN(_02590_ ) );
NOR2_X1 _09737_ ( .A1(_02589_ ), .A2(_02590_ ), .ZN(_02591_ ) );
AND3_X1 _09738_ ( .A1(_02588_ ), .A2(_01675_ ), .A3(_02591_ ), .ZN(_02592_ ) );
INV_X1 _09739_ ( .A(\u_lsu.u_clint.mtime[3] ), .ZN(_02593_ ) );
NAND4_X1 _09740_ ( .A1(_01276_ ), .A2(_01258_ ), .A3(\io_master_araddr[3] ), .A4(_02593_ ), .ZN(_02594_ ) );
OAI211_X1 _09741_ ( .A(_01595_ ), .B(_02594_ ), .C1(\u_lsu.u_clint.mtime[35] ), .C2(_01599_ ), .ZN(_02595_ ) );
AOI21_X1 _09742_ ( .A(_01664_ ), .B1(io_master_rready ), .B2(\io_master_rdata[3] ), .ZN(_02596_ ) );
AND2_X1 _09743_ ( .A1(_02595_ ), .A2(_02596_ ), .ZN(_02597_ ) );
NOR3_X1 _09744_ ( .A1(_02592_ ), .A2(_02412_ ), .A3(_02597_ ), .ZN(_02598_ ) );
MUX2_X1 _09745_ ( .A(_02587_ ), .B(_02598_ ), .S(fanout_net_12 ), .Z(\ar_data[3] ) );
NAND2_X1 _09746_ ( .A1(\ar_data[3] ), .A2(_01531_ ), .ZN(_02599_ ) );
AOI22_X1 _09747_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02600_ ) );
AOI22_X1 _09748_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02601_ ) );
NAND3_X1 _09749_ ( .A1(_02600_ ), .A2(_02601_ ), .A3(_01841_ ), .ZN(_02602_ ) );
AOI22_X1 _09750_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02603_ ) );
AOI22_X1 _09751_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02604_ ) );
NAND3_X1 _09752_ ( .A1(_02603_ ), .A2(_02604_ ), .A3(_01829_ ), .ZN(_02605_ ) );
NAND3_X1 _09753_ ( .A1(_02602_ ), .A2(_02605_ ), .A3(_01855_ ), .ZN(_02606_ ) );
OAI211_X1 _09754_ ( .A(fanout_net_21 ), .B(_01838_ ), .C1(_01903_ ), .C2(\u_reg.rf[1][3] ), .ZN(_02607_ ) );
OAI21_X1 _09755_ ( .A(_02607_ ), .B1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01833_ ), .ZN(_02608_ ) );
NAND3_X1 _09756_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_02609_ ) );
AND3_X1 _09757_ ( .A1(_02608_ ), .A2(_01841_ ), .A3(_02609_ ), .ZN(_02610_ ) );
AOI22_X1 _09758_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01826_ ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02611_ ) );
NAND3_X1 _09759_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_02612_ ) );
NAND3_X1 _09760_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01833_ ), .ZN(_02613_ ) );
NAND4_X1 _09761_ ( .A1(_02611_ ), .A2(_01901_ ), .A3(_02612_ ), .A4(_02613_ ), .ZN(_02614_ ) );
NAND2_X1 _09762_ ( .A1(_02614_ ), .A2(_01836_ ), .ZN(_02615_ ) );
OAI211_X1 _09763_ ( .A(_01823_ ), .B(_02606_ ), .C1(_02610_ ), .C2(_02615_ ), .ZN(_02616_ ) );
AOI21_X1 _09764_ ( .A(_01999_ ), .B1(_02599_ ), .B2(_02616_ ), .ZN(_02617_ ) );
AND2_X1 _09765_ ( .A1(_02617_ ), .A2(_01533_ ), .ZN(_02618_ ) );
OAI211_X1 _09766_ ( .A(_01622_ ), .B(\u_csr.csr[3][0] ), .C1(_01620_ ), .C2(_00858_ ), .ZN(_02619_ ) );
NOR3_X1 _09767_ ( .A1(_02619_ ), .A2(_01624_ ), .A3(_01625_ ), .ZN(_02620_ ) );
NOR2_X1 _09768_ ( .A1(_01544_ ), .A2(_01627_ ), .ZN(_02621_ ) );
INV_X1 _09769_ ( .A(_02621_ ), .ZN(_02622_ ) );
AOI211_X1 _09770_ ( .A(_02620_ ), .B(_02622_ ), .C1(\u_csr.csr[1][3] ), .C2(_01631_ ), .ZN(_02623_ ) );
NAND4_X1 _09771_ ( .A1(_01928_ ), .A2(\u_csr.csr[2][3] ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_02624_ ) );
NAND3_X1 _09772_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][3] ), .A3(_01874_ ), .ZN(_02625_ ) );
AND2_X1 _09773_ ( .A1(_02624_ ), .A2(_02625_ ), .ZN(_02626_ ) );
AOI21_X1 _09774_ ( .A(_01619_ ), .B1(_02623_ ), .B2(_02626_ ), .ZN(_02627_ ) );
NAND2_X1 _09775_ ( .A1(_00829_ ), .A2(_00830_ ), .ZN(_02628_ ) );
NOR3_X1 _09776_ ( .A1(_01393_ ), .A2(_01413_ ), .A3(_01401_ ), .ZN(_02629_ ) );
AND4_X1 _09777_ ( .A1(_02628_ ), .A2(_02629_ ), .A3(_01425_ ), .A4(_01406_ ), .ZN(_02630_ ) );
NOR2_X1 _09778_ ( .A1(_02627_ ), .A2(_02630_ ), .ZN(_02631_ ) );
INV_X1 _09779_ ( .A(\de_pc[3] ), .ZN(_02632_ ) );
OAI22_X1 _09780_ ( .A1(_02631_ ), .A2(_01353_ ), .B1(_02632_ ), .B2(_01453_ ), .ZN(_02633_ ) );
OAI21_X1 _09781_ ( .A(_01720_ ), .B1(_02618_ ), .B2(_02633_ ), .ZN(_02634_ ) );
NAND2_X1 _09782_ ( .A1(_02617_ ), .A2(_01557_ ), .ZN(_02635_ ) );
AOI21_X1 _09783_ ( .A(_00944_ ), .B1(_00728_ ), .B2(_00693_ ), .ZN(_02636_ ) );
AOI21_X1 _09784_ ( .A(_00893_ ), .B1(_02579_ ), .B2(_00924_ ), .ZN(_02637_ ) );
NOR2_X1 _09785_ ( .A1(_02636_ ), .A2(_02637_ ), .ZN(_02638_ ) );
INV_X1 _09786_ ( .A(_02638_ ), .ZN(_02639_ ) );
NAND3_X1 _09787_ ( .A1(_02578_ ), .A2(_02407_ ), .A3(_02639_ ), .ZN(_02640_ ) );
NAND3_X1 _09788_ ( .A1(_02578_ ), .A2(\de_pc[3] ), .A3(_01861_ ), .ZN(_02641_ ) );
AND3_X1 _09789_ ( .A1(_02635_ ), .A2(_02640_ ), .A3(_02641_ ), .ZN(_02642_ ) );
OAI21_X1 _09790_ ( .A(_02634_ ), .B1(_02642_ ), .B2(_01806_ ), .ZN(_00150_ ) );
AOI22_X1 _09791_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01826_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02643_ ) );
AOI22_X1 _09792_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02644_ ) );
NAND3_X1 _09793_ ( .A1(_02643_ ), .A2(_02644_ ), .A3(_01841_ ), .ZN(_02645_ ) );
AOI22_X1 _09794_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02646_ ) );
AOI22_X1 _09795_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02647_ ) );
NAND3_X1 _09796_ ( .A1(_02646_ ), .A2(_02647_ ), .A3(_01829_ ), .ZN(_02648_ ) );
NAND3_X1 _09797_ ( .A1(_02645_ ), .A2(_02648_ ), .A3(_01855_ ), .ZN(_02649_ ) );
OAI211_X1 _09798_ ( .A(fanout_net_21 ), .B(_01838_ ), .C1(_01903_ ), .C2(\u_reg.rf[1][2] ), .ZN(_02650_ ) );
OAI21_X1 _09799_ ( .A(_02650_ ), .B1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01833_ ), .ZN(_02651_ ) );
NAND3_X1 _09800_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_02652_ ) );
AND3_X1 _09801_ ( .A1(_02651_ ), .A2(_01841_ ), .A3(_02652_ ), .ZN(_02653_ ) );
AOI22_X1 _09802_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01826_ ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02654_ ) );
NAND3_X1 _09803_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_02655_ ) );
NAND3_X1 _09804_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01833_ ), .ZN(_02656_ ) );
NAND4_X1 _09805_ ( .A1(_02654_ ), .A2(_01829_ ), .A3(_02655_ ), .A4(_02656_ ), .ZN(_02657_ ) );
NAND2_X1 _09806_ ( .A1(_02657_ ), .A2(_01836_ ), .ZN(_02658_ ) );
OAI211_X1 _09807_ ( .A(_01823_ ), .B(_02649_ ), .C1(_02653_ ), .C2(_02658_ ), .ZN(_02659_ ) );
MUX2_X1 _09808_ ( .A(\ea_addr[2] ), .B(\u_exu.ecsr[2] ), .S(_01527_ ), .Z(_02660_ ) );
NOR2_X1 _09809_ ( .A1(_02298_ ), .A2(_01285_ ), .ZN(_02661_ ) );
INV_X1 _09810_ ( .A(_02661_ ), .ZN(_02662_ ) );
AND3_X1 _09811_ ( .A1(_01815_ ), .A2(_01281_ ), .A3(_01819_ ), .ZN(_02663_ ) );
AOI21_X1 _09812_ ( .A(_02663_ ), .B1(_01255_ ), .B2(_01814_ ), .ZN(_02664_ ) );
AND3_X1 _09813_ ( .A1(_02662_ ), .A2(_02664_ ), .A3(_01664_ ), .ZN(_02665_ ) );
INV_X1 _09814_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_28_A_$_ANDNOT__Y_B ), .ZN(_02666_ ) );
NOR2_X1 _09815_ ( .A1(_01598_ ), .A2(_02666_ ), .ZN(_02667_ ) );
INV_X1 _09816_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ), .ZN(_02668_ ) );
NOR3_X1 _09817_ ( .A1(_01518_ ), .A2(\u_arbiter.raddr[2] ), .A3(_02668_ ), .ZN(_02669_ ) );
NOR4_X1 _09818_ ( .A1(_01601_ ), .A2(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .A3(_02667_ ), .A4(_02669_ ), .ZN(_02670_ ) );
AOI21_X1 _09819_ ( .A(_02670_ ), .B1(io_master_rready ), .B2(\io_master_rdata[2] ), .ZN(_02671_ ) );
AND2_X1 _09820_ ( .A1(_02671_ ), .A2(_01276_ ), .ZN(_02672_ ) );
NOR3_X1 _09821_ ( .A1(_02665_ ), .A2(_02412_ ), .A3(_02672_ ), .ZN(_02673_ ) );
MUX2_X1 _09822_ ( .A(_02660_ ), .B(_02673_ ), .S(fanout_net_12 ), .Z(\ar_data[2] ) );
NAND2_X1 _09823_ ( .A1(\ar_data[2] ), .A2(_01531_ ), .ZN(_02674_ ) );
AOI21_X1 _09824_ ( .A(_01999_ ), .B1(_02659_ ), .B2(_02674_ ), .ZN(_02675_ ) );
AND2_X1 _09825_ ( .A1(_02675_ ), .A2(_01533_ ), .ZN(_02676_ ) );
AOI211_X1 _09826_ ( .A(_01419_ ), .B(_01424_ ), .C1(_00831_ ), .C2(_00832_ ), .ZN(_02677_ ) );
NAND3_X1 _09827_ ( .A1(_01778_ ), .A2(\u_csr.csr[1][2] ), .A3(_01779_ ), .ZN(_02678_ ) );
AND3_X1 _09828_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][2] ), .A3(_01435_ ), .ZN(_02679_ ) );
AOI21_X1 _09829_ ( .A(_02679_ ), .B1(_01783_ ), .B2(_01626_ ), .ZN(_02680_ ) );
NAND4_X1 _09830_ ( .A1(_01431_ ), .A2(\u_csr.csr[2][2] ), .A3(_01785_ ), .A4(_01786_ ), .ZN(_02681_ ) );
NAND3_X1 _09831_ ( .A1(_02678_ ), .A2(_02680_ ), .A3(_02681_ ), .ZN(_02682_ ) );
AND3_X1 _09832_ ( .A1(_01776_ ), .A2(_01425_ ), .A3(_02682_ ), .ZN(_02683_ ) );
NOR2_X1 _09833_ ( .A1(_02677_ ), .A2(_02683_ ), .ZN(_02684_ ) );
INV_X1 _09834_ ( .A(\de_pc[2] ), .ZN(_02685_ ) );
OAI22_X1 _09835_ ( .A1(_02684_ ), .A2(_01353_ ), .B1(_02685_ ), .B2(_01453_ ), .ZN(_02686_ ) );
OAI21_X1 _09836_ ( .A(_01720_ ), .B1(_02676_ ), .B2(_02686_ ), .ZN(_02687_ ) );
NAND2_X1 _09837_ ( .A1(_02675_ ), .A2(_01557_ ), .ZN(_02688_ ) );
INV_X1 _09838_ ( .A(_01469_ ), .ZN(_02689_ ) );
AND2_X1 _09839_ ( .A1(_02689_ ), .A2(\u_idu.imm_branch[2] ), .ZN(_02690_ ) );
AOI21_X1 _09840_ ( .A(_00894_ ), .B1(_02579_ ), .B2(_00924_ ), .ZN(_02691_ ) );
NOR2_X1 _09841_ ( .A1(_02690_ ), .A2(_02691_ ), .ZN(_02692_ ) );
INV_X1 _09842_ ( .A(_02692_ ), .ZN(_02693_ ) );
NAND3_X1 _09843_ ( .A1(_02578_ ), .A2(_02407_ ), .A3(_02693_ ), .ZN(_02694_ ) );
NAND3_X1 _09844_ ( .A1(_02578_ ), .A2(\de_pc[2] ), .A3(_01566_ ), .ZN(_02695_ ) );
AND3_X1 _09845_ ( .A1(_02688_ ), .A2(_02694_ ), .A3(_02695_ ), .ZN(_02696_ ) );
OAI21_X1 _09846_ ( .A(_02687_ ), .B1(_02696_ ), .B2(_01806_ ), .ZN(_00151_ ) );
AND3_X1 _09847_ ( .A1(_02160_ ), .A2(_01523_ ), .A3(\io_master_arsize[1] ), .ZN(_02697_ ) );
NOR3_X1 _09848_ ( .A1(_01275_ ), .A2(_01295_ ), .A3(_02697_ ), .ZN(_02698_ ) );
NAND2_X1 _09849_ ( .A1(_02698_ ), .A2(fanout_net_12 ), .ZN(_02699_ ) );
MUX2_X1 _09850_ ( .A(\ea_addr[28] ), .B(\u_exu.ecsr[28] ), .S(_01299_ ), .Z(_02700_ ) );
OR2_X1 _09851_ ( .A1(_02700_ ), .A2(fanout_net_12 ), .ZN(_02701_ ) );
AOI21_X1 _09852_ ( .A(_01245_ ), .B1(_02699_ ), .B2(_02701_ ), .ZN(_02702_ ) );
AOI22_X1 _09853_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02703_ ) );
AOI22_X1 _09854_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02704_ ) );
NAND3_X1 _09855_ ( .A1(_02703_ ), .A2(_02704_ ), .A3(_01312_ ), .ZN(_02705_ ) );
AOI22_X1 _09856_ ( .A1(_01005_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02706_ ) );
AOI22_X1 _09857_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02707_ ) );
NAND3_X1 _09858_ ( .A1(_02706_ ), .A2(_02707_ ), .A3(_00915_ ), .ZN(_02708_ ) );
AND3_X1 _09859_ ( .A1(_02705_ ), .A2(_02708_ ), .A3(_01320_ ), .ZN(_02709_ ) );
NAND3_X1 _09860_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01339_ ), .ZN(_02710_ ) );
INV_X1 _09861_ ( .A(\u_reg.rf[1][28] ), .ZN(_02711_ ) );
AOI21_X1 _09862_ ( .A(_01506_ ), .B1(_01589_ ), .B2(_02711_ ), .ZN(_02712_ ) );
NOR2_X1 _09863_ ( .A1(_01589_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02713_ ) );
OAI211_X1 _09864_ ( .A(_01580_ ), .B(_02710_ ), .C1(_02712_ ), .C2(_02713_ ), .ZN(_02714_ ) );
AOI22_X1 _09865_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02715_ ) );
AOI22_X1 _09866_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02716_ ) );
NAND3_X1 _09867_ ( .A1(_02715_ ), .A2(_02716_ ), .A3(_01484_ ), .ZN(_02717_ ) );
AND2_X1 _09868_ ( .A1(_02717_ ), .A2(_01046_ ), .ZN(_02718_ ) );
AOI21_X1 _09869_ ( .A(_02709_ ), .B1(_02714_ ), .B2(_02718_ ), .ZN(_02719_ ) );
OAI21_X1 _09870_ ( .A(_00736_ ), .B1(_01304_ ), .B2(_02719_ ), .ZN(_02720_ ) );
OR3_X1 _09871_ ( .A1(_02702_ ), .A2(_00723_ ), .A3(_02720_ ), .ZN(_02721_ ) );
NAND4_X1 _09872_ ( .A1(_01415_ ), .A2(_00838_ ), .A3(_00837_ ), .A4(_01421_ ), .ZN(_02722_ ) );
AND3_X1 _09873_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][28] ), .A3(_01435_ ), .ZN(_02723_ ) );
AOI21_X1 _09874_ ( .A(_02723_ ), .B1(_01539_ ), .B2(_01783_ ), .ZN(_02724_ ) );
NAND3_X1 _09875_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][28] ), .A3(_02210_ ), .ZN(_02725_ ) );
NAND4_X1 _09876_ ( .A1(_02210_ ), .A2(\u_csr.csr[2][28] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_02726_ ) );
NAND3_X1 _09877_ ( .A1(_02724_ ), .A2(_02725_ ), .A3(_02726_ ), .ZN(_02727_ ) );
NAND3_X1 _09878_ ( .A1(_01775_ ), .A2(_01538_ ), .A3(_02727_ ), .ZN(_02728_ ) );
AOI21_X1 _09879_ ( .A(_01535_ ), .B1(_02722_ ), .B2(_02728_ ), .ZN(_02729_ ) );
AOI221_X4 _09880_ ( .A(_02729_ ), .B1(\de_pc[28] ), .B2(_01454_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_02730_ ) );
OR3_X1 _09881_ ( .A1(_02702_ ), .A2(_01460_ ), .A3(_02720_ ), .ZN(_02731_ ) );
AOI21_X1 _09882_ ( .A(_01562_ ), .B1(\u_idu.imm_auipc_lui[28] ), .B2(_01563_ ), .ZN(_02732_ ) );
NOR3_X1 _09883_ ( .A1(_02732_ ), .A2(_01555_ ), .A3(_01566_ ), .ZN(_02733_ ) );
AOI211_X1 _09884_ ( .A(_02733_ ), .B(_01053_ ), .C1(\de_pc[28] ), .C2(_01464_ ), .ZN(_02734_ ) );
AOI221_X1 _09885_ ( .A(_01644_ ), .B1(_02721_ ), .B2(_02730_ ), .C1(_02731_ ), .C2(_02734_ ), .ZN(_00152_ ) );
MUX2_X1 _09886_ ( .A(\ea_addr[1] ), .B(\u_exu.ecsr[1] ), .S(_01299_ ), .Z(_02735_ ) );
OAI22_X1 _09887_ ( .A1(_01894_ ), .A2(_01256_ ), .B1(_01884_ ), .B2(_02324_ ), .ZN(_02736_ ) );
AOI21_X1 _09888_ ( .A(_01282_ ), .B1(_01887_ ), .B2(_01888_ ), .ZN(_02737_ ) );
NOR3_X1 _09889_ ( .A1(_02736_ ), .A2(_01523_ ), .A3(_02737_ ), .ZN(_02738_ ) );
OR3_X1 _09890_ ( .A1(_01946_ ), .A2(\u_arbiter.raddr[2] ), .A3(\u_lsu.u_clint.mtime[1] ), .ZN(_02739_ ) );
OAI211_X1 _09891_ ( .A(_01595_ ), .B(_02739_ ), .C1(\u_lsu.u_clint.mtime[33] ), .C2(_01599_ ), .ZN(_02740_ ) );
AOI21_X1 _09892_ ( .A(_01664_ ), .B1(io_master_rready ), .B2(\io_master_rdata[1] ), .ZN(_02741_ ) );
AND2_X1 _09893_ ( .A1(_02740_ ), .A2(_02741_ ), .ZN(_02742_ ) );
NOR3_X1 _09894_ ( .A1(_02738_ ), .A2(_02412_ ), .A3(_02742_ ), .ZN(_02743_ ) );
MUX2_X1 _09895_ ( .A(_02735_ ), .B(_02743_ ), .S(fanout_net_12 ), .Z(\ar_data[1] ) );
NAND2_X1 _09896_ ( .A1(\ar_data[1] ), .A2(_01531_ ), .ZN(_02744_ ) );
AOI22_X1 _09897_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02745_ ) );
AOI22_X1 _09898_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02746_ ) );
NAND3_X1 _09899_ ( .A1(_02745_ ), .A2(_02746_ ), .A3(_01841_ ), .ZN(_02747_ ) );
AOI22_X1 _09900_ ( .A1(_01917_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02748_ ) );
AOI22_X1 _09901_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02749_ ) );
NAND3_X1 _09902_ ( .A1(_02748_ ), .A2(_02749_ ), .A3(_01901_ ), .ZN(_02750_ ) );
NAND3_X1 _09903_ ( .A1(_02747_ ), .A2(_02750_ ), .A3(_01855_ ), .ZN(_02751_ ) );
AOI22_X1 _09904_ ( .A1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01826_ ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02752_ ) );
NAND3_X1 _09905_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_02753_ ) );
NAND3_X1 _09906_ ( .A1(_01902_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01833_ ), .ZN(_02754_ ) );
AND4_X1 _09907_ ( .A1(_01829_ ), .A2(_02752_ ), .A3(_02753_ ), .A4(_02754_ ), .ZN(_02755_ ) );
OAI21_X1 _09908_ ( .A(_01506_ ), .B1(_01342_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02756_ ) );
OAI21_X1 _09909_ ( .A(_02756_ ), .B1(\u_reg.rf[1][1] ), .B2(_01587_ ), .ZN(_02757_ ) );
AOI211_X1 _09910_ ( .A(_01585_ ), .B(_02757_ ), .C1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_01914_ ), .ZN(_02758_ ) );
OR2_X1 _09911_ ( .A1(_02758_ ), .A2(_01756_ ), .ZN(_02759_ ) );
OAI211_X1 _09912_ ( .A(_01823_ ), .B(_02751_ ), .C1(_02755_ ), .C2(_02759_ ), .ZN(_02760_ ) );
AOI21_X1 _09913_ ( .A(_01999_ ), .B1(_02744_ ), .B2(_02760_ ), .ZN(_02761_ ) );
AND2_X1 _09914_ ( .A1(_02761_ ), .A2(_01533_ ), .ZN(_02762_ ) );
AND3_X1 _09915_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][1] ), .A3(_01874_ ), .ZN(_02763_ ) );
AOI21_X1 _09916_ ( .A(_02763_ ), .B1(_01631_ ), .B2(\u_csr.csr[1][1] ), .ZN(_02764_ ) );
AND4_X1 _09917_ ( .A1(\u_csr.csr[2][1] ), .A2(_01928_ ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_02765_ ) );
NOR3_X1 _09918_ ( .A1(_02765_ ), .A2(_02620_ ), .A3(_01627_ ), .ZN(_02766_ ) );
AOI21_X1 _09919_ ( .A(_01619_ ), .B1(_02764_ ), .B2(_02766_ ), .ZN(_02767_ ) );
AOI211_X1 _09920_ ( .A(_01419_ ), .B(_01424_ ), .C1(_00833_ ), .C2(_00834_ ), .ZN(_02768_ ) );
NOR2_X1 _09921_ ( .A1(_02767_ ), .A2(_02768_ ), .ZN(_02769_ ) );
INV_X1 _09922_ ( .A(\de_pc[1] ), .ZN(_02770_ ) );
OAI22_X1 _09923_ ( .A1(_02769_ ), .A2(_01353_ ), .B1(_02770_ ), .B2(_01453_ ), .ZN(_02771_ ) );
OAI21_X1 _09924_ ( .A(_01720_ ), .B1(_02762_ ), .B2(_02771_ ), .ZN(_02772_ ) );
NAND2_X1 _09925_ ( .A1(_02761_ ), .A2(_01557_ ), .ZN(_02773_ ) );
OR2_X1 _09926_ ( .A1(_02580_ ), .A2(_01641_ ), .ZN(_02774_ ) );
OAI21_X1 _09927_ ( .A(\u_idu.imm_branch[1] ), .B1(_00727_ ), .B2(_00692_ ), .ZN(_02775_ ) );
NAND2_X1 _09928_ ( .A1(_02774_ ), .A2(_02775_ ), .ZN(_02776_ ) );
NAND3_X1 _09929_ ( .A1(_02578_ ), .A2(_02407_ ), .A3(_02776_ ), .ZN(_02777_ ) );
NAND3_X1 _09930_ ( .A1(_02578_ ), .A2(\de_pc[1] ), .A3(_01566_ ), .ZN(_02778_ ) );
AND3_X1 _09931_ ( .A1(_02773_ ), .A2(_02777_ ), .A3(_02778_ ), .ZN(_02779_ ) );
OAI21_X1 _09932_ ( .A(_02772_ ), .B1(_02779_ ), .B2(_01805_ ), .ZN(_00153_ ) );
OAI21_X1 _09933_ ( .A(_01506_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02780_ ) );
OAI21_X1 _09934_ ( .A(_02780_ ), .B1(\u_reg.rf[1][0] ), .B2(_01903_ ), .ZN(_02781_ ) );
AND4_X1 _09935_ ( .A1(fanout_net_21 ), .A2(_01339_ ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A4(_01837_ ), .ZN(_02782_ ) );
OR3_X1 _09936_ ( .A1(_02781_ ), .A2(_01744_ ), .A3(_02782_ ), .ZN(_02783_ ) );
AOI22_X1 _09937_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01826_ ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02784_ ) );
NAND3_X1 _09938_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01831_ ), .ZN(_02785_ ) );
NAND3_X1 _09939_ ( .A1(_01830_ ), .A2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01833_ ), .ZN(_02786_ ) );
NAND4_X1 _09940_ ( .A1(_02784_ ), .A2(_01829_ ), .A3(_02785_ ), .A4(_02786_ ), .ZN(_02787_ ) );
NAND3_X1 _09941_ ( .A1(_02783_ ), .A2(_01836_ ), .A3(_02787_ ), .ZN(_02788_ ) );
AOI22_X1 _09942_ ( .A1(_01845_ ), .A2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01826_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02789_ ) );
AOI22_X1 _09943_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01827_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02790_ ) );
AOI21_X1 _09944_ ( .A(_01829_ ), .B1(_02789_ ), .B2(_02790_ ), .ZN(_02791_ ) );
AOI22_X1 _09945_ ( .A1(_01847_ ), .A2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01850_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02792_ ) );
AOI22_X1 _09946_ ( .A1(_01914_ ), .A2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01852_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02793_ ) );
AOI21_X1 _09947_ ( .A(_01910_ ), .B1(_02792_ ), .B2(_02793_ ), .ZN(_02794_ ) );
OAI21_X1 _09948_ ( .A(_01855_ ), .B1(_02791_ ), .B2(_02794_ ), .ZN(_02795_ ) );
NAND3_X1 _09949_ ( .A1(_01823_ ), .A2(_02788_ ), .A3(_02795_ ), .ZN(_02796_ ) );
NAND3_X1 _09950_ ( .A1(_01945_ ), .A2(_01255_ ), .A3(_01951_ ), .ZN(_02797_ ) );
OAI221_X1 _09951_ ( .A(_02797_ ), .B1(_01884_ ), .B2(_02373_ ), .C1(_01960_ ), .C2(_01282_ ), .ZN(_02798_ ) );
NAND4_X1 _09952_ ( .A1(_01523_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D[0] ), .A3(\io_master_araddr[3] ), .A4(_01258_ ), .ZN(_02799_ ) );
INV_X1 _09953_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A ), .ZN(_02800_ ) );
OAI211_X1 _09954_ ( .A(_01595_ ), .B(_02799_ ), .C1(_02800_ ), .C2(_01599_ ), .ZN(_02801_ ) );
NAND2_X1 _09955_ ( .A1(io_master_rready ), .A2(\io_master_rdata[0] ), .ZN(_02802_ ) );
AOI21_X1 _09956_ ( .A(_01675_ ), .B1(_02801_ ), .B2(_02802_ ), .ZN(_02803_ ) );
OAI21_X1 _09957_ ( .A(_02465_ ), .B1(_02798_ ), .B2(_02803_ ), .ZN(_02804_ ) );
NAND2_X1 _09958_ ( .A1(_02804_ ), .A2(fanout_net_12 ), .ZN(_02805_ ) );
MUX2_X1 _09959_ ( .A(\ea_addr[0] ), .B(\u_exu.ecsr[0] ), .S(_01299_ ), .Z(_02806_ ) );
OR2_X1 _09960_ ( .A1(_02806_ ), .A2(fanout_net_12 ), .ZN(_02807_ ) );
NAND4_X1 _09961_ ( .A1(_02805_ ), .A2(_01223_ ), .A3(_01243_ ), .A4(_02807_ ), .ZN(_02808_ ) );
AOI21_X1 _09962_ ( .A(_01999_ ), .B1(_02796_ ), .B2(_02808_ ), .ZN(_02809_ ) );
AND2_X1 _09963_ ( .A1(_02809_ ), .A2(_01533_ ), .ZN(_02810_ ) );
AND3_X1 _09964_ ( .A1(_01873_ ), .A2(\u_csr.csr[0][0] ), .A3(_01874_ ), .ZN(_02811_ ) );
AOI21_X1 _09965_ ( .A(_02811_ ), .B1(_01631_ ), .B2(\u_csr.csr[1][0] ), .ZN(_02812_ ) );
AND4_X1 _09966_ ( .A1(\u_csr.csr[2][0] ), .A2(_01928_ ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_02813_ ) );
NOR3_X1 _09967_ ( .A1(_02813_ ), .A2(_02620_ ), .A3(_01627_ ), .ZN(_02814_ ) );
AOI21_X1 _09968_ ( .A(_01619_ ), .B1(_02812_ ), .B2(_02814_ ), .ZN(_02815_ ) );
AOI211_X1 _09969_ ( .A(_01419_ ), .B(_01424_ ), .C1(_00835_ ), .C2(_00836_ ), .ZN(_02816_ ) );
NOR2_X1 _09970_ ( .A1(_02815_ ), .A2(_02816_ ), .ZN(_02817_ ) );
INV_X1 _09971_ ( .A(\de_pc[0] ), .ZN(_02818_ ) );
OAI22_X1 _09972_ ( .A1(_02817_ ), .A2(_01353_ ), .B1(_02818_ ), .B2(_01453_ ), .ZN(_02819_ ) );
OAI21_X1 _09973_ ( .A(_01720_ ), .B1(_02810_ ), .B2(_02819_ ), .ZN(_02820_ ) );
NAND2_X1 _09974_ ( .A1(_02809_ ), .A2(_01557_ ), .ZN(_02821_ ) );
AND4_X1 _09975_ ( .A1(fanout_net_22 ), .A2(_00687_ ), .A3(_00691_ ), .A4(_00719_ ), .ZN(_02822_ ) );
AOI21_X1 _09976_ ( .A(_02822_ ), .B1(_00882_ ), .B2(_00734_ ), .ZN(_02823_ ) );
INV_X1 _09977_ ( .A(_02823_ ), .ZN(_02824_ ) );
AND3_X1 _09978_ ( .A1(_00726_ ), .A2(\u_idu.imm_branch[11] ), .A3(\u_idu.inst[5] ), .ZN(_02825_ ) );
AND3_X1 _09979_ ( .A1(_00665_ ), .A2(fanout_net_22 ), .A3(_00670_ ), .ZN(_02826_ ) );
NOR3_X1 _09980_ ( .A1(_02824_ ), .A2(_02825_ ), .A3(_02826_ ), .ZN(_02827_ ) );
INV_X1 _09981_ ( .A(_02827_ ), .ZN(_02828_ ) );
NAND3_X1 _09982_ ( .A1(_02578_ ), .A2(_02407_ ), .A3(_02828_ ), .ZN(_02829_ ) );
NAND3_X1 _09983_ ( .A1(_02578_ ), .A2(\de_pc[0] ), .A3(_01566_ ), .ZN(_02830_ ) );
AND3_X1 _09984_ ( .A1(_02821_ ), .A2(_02829_ ), .A3(_02830_ ), .ZN(_02831_ ) );
OAI21_X1 _09985_ ( .A(_02820_ ), .B1(_02831_ ), .B2(_01805_ ), .ZN(_00154_ ) );
AOI22_X1 _09986_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02832_ ) );
AOI22_X1 _09987_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02833_ ) );
NAND3_X1 _09988_ ( .A1(_02832_ ), .A2(_02833_ ), .A3(_01312_ ), .ZN(_02834_ ) );
AOI22_X1 _09989_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02835_ ) );
AOI22_X1 _09990_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02836_ ) );
NAND3_X1 _09991_ ( .A1(_02835_ ), .A2(_02836_ ), .A3(_01318_ ), .ZN(_02837_ ) );
AND3_X1 _09992_ ( .A1(_02834_ ), .A2(_02837_ ), .A3(_01320_ ), .ZN(_02838_ ) );
OAI211_X1 _09993_ ( .A(fanout_net_21 ), .B(_01322_ ), .C1(_01323_ ), .C2(\u_reg.rf[1][27] ), .ZN(_02839_ ) );
OAI21_X1 _09994_ ( .A(_02839_ ), .B1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01342_ ), .ZN(_02840_ ) );
NAND4_X1 _09995_ ( .A1(_01328_ ), .A2(fanout_net_21 ), .A3(_01322_ ), .A4(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02841_ ) );
NAND3_X1 _09996_ ( .A1(_02840_ ), .A2(_01580_ ), .A3(_02841_ ), .ZN(_02842_ ) );
AND2_X1 _09997_ ( .A1(_02842_ ), .A2(_01504_ ), .ZN(_02843_ ) );
AOI22_X1 _09998_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01333_ ), .B1(_01334_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02844_ ) );
NAND3_X1 _09999_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01587_ ), .ZN(_02845_ ) );
NAND3_X1 _10000_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01589_ ), .ZN(_02846_ ) );
NAND4_X1 _10001_ ( .A1(_02844_ ), .A2(_01585_ ), .A3(_02845_ ), .A4(_02846_ ), .ZN(_02847_ ) );
AOI21_X1 _10002_ ( .A(_02838_ ), .B1(_02843_ ), .B2(_02847_ ), .ZN(_02848_ ) );
OAI21_X1 _10003_ ( .A(_01303_ ), .B1(_01482_ ), .B2(_02848_ ), .ZN(_02849_ ) );
AOI21_X1 _10004_ ( .A(_01279_ ), .B1(_01732_ ), .B2(_01733_ ), .ZN(_02850_ ) );
NOR3_X1 _10005_ ( .A1(_01275_ ), .A2(_01294_ ), .A3(_02850_ ), .ZN(_02851_ ) );
NAND2_X1 _10006_ ( .A1(_02851_ ), .A2(fanout_net_12 ), .ZN(_02852_ ) );
MUX2_X1 _10007_ ( .A(\ea_addr[27] ), .B(\u_exu.ecsr[27] ), .S(_01527_ ), .Z(_02853_ ) );
OR2_X1 _10008_ ( .A1(_02853_ ), .A2(fanout_net_12 ), .ZN(_02854_ ) );
AND2_X1 _10009_ ( .A1(_02852_ ), .A2(_02854_ ), .ZN(\ar_data[27] ) );
INV_X1 _10010_ ( .A(\ar_data[27] ), .ZN(_02855_ ) );
AOI21_X1 _10011_ ( .A(_02849_ ), .B1(_02855_ ), .B2(_01531_ ), .ZN(_02856_ ) );
NAND2_X1 _10012_ ( .A1(_02856_ ), .A2(_00743_ ), .ZN(_02857_ ) );
NAND4_X1 _10013_ ( .A1(_01416_ ), .A2(_00841_ ), .A3(_00839_ ), .A4(_01421_ ), .ZN(_02858_ ) );
AND3_X1 _10014_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][27] ), .A3(_01435_ ), .ZN(_02859_ ) );
AOI21_X1 _10015_ ( .A(_02859_ ), .B1(_01928_ ), .B2(_01783_ ), .ZN(_02860_ ) );
NAND3_X1 _10016_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][27] ), .A3(_01431_ ), .ZN(_02861_ ) );
NAND4_X1 _10017_ ( .A1(_02210_ ), .A2(\u_csr.csr[2][27] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_02862_ ) );
NAND3_X1 _10018_ ( .A1(_02860_ ), .A2(_02861_ ), .A3(_02862_ ), .ZN(_02863_ ) );
NAND3_X1 _10019_ ( .A1(_01776_ ), .A2(_01538_ ), .A3(_02863_ ), .ZN(_02864_ ) );
AOI21_X1 _10020_ ( .A(_01535_ ), .B1(_02858_ ), .B2(_02864_ ), .ZN(_02865_ ) );
AOI221_X4 _10021_ ( .A(_02865_ ), .B1(\de_pc[27] ), .B2(_01454_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_02866_ ) );
NAND2_X1 _10022_ ( .A1(_02856_ ), .A2(_01556_ ), .ZN(_02867_ ) );
AOI21_X1 _10023_ ( .A(_01562_ ), .B1(\u_idu.imm_auipc_lui[27] ), .B2(_01563_ ), .ZN(_02868_ ) );
NOR3_X1 _10024_ ( .A1(_02868_ ), .A2(_01555_ ), .A3(_01566_ ), .ZN(_02869_ ) );
AOI211_X1 _10025_ ( .A(_02869_ ), .B(_01053_ ), .C1(\de_pc[27] ), .C2(_01464_ ), .ZN(_02870_ ) );
AOI221_X4 _10026_ ( .A(_01644_ ), .B1(_02857_ ), .B2(_02866_ ), .C1(_02867_ ), .C2(_02870_ ), .ZN(_00155_ ) );
AOI22_X1 _10027_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01486_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02871_ ) );
AOI22_X1 _10028_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02872_ ) );
AOI21_X1 _10029_ ( .A(_01484_ ), .B1(_02871_ ), .B2(_02872_ ), .ZN(_02873_ ) );
AOI22_X1 _10030_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02874_ ) );
AOI22_X1 _10031_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02875_ ) );
AOI21_X1 _10032_ ( .A(_01327_ ), .B1(_02874_ ), .B2(_02875_ ), .ZN(_02876_ ) );
OAI21_X1 _10033_ ( .A(_01483_ ), .B1(_02873_ ), .B2(_02876_ ), .ZN(_02877_ ) );
AOI22_X1 _10034_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01486_ ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02878_ ) );
NAND3_X1 _10035_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01328_ ), .ZN(_02879_ ) );
NAND3_X1 _10036_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01325_ ), .ZN(_02880_ ) );
NAND4_X1 _10037_ ( .A1(_02878_ ), .A2(_01336_ ), .A3(_02879_ ), .A4(_02880_ ), .ZN(_02881_ ) );
OAI211_X1 _10038_ ( .A(\u_idu.imm_auipc_lui[15] ), .B(_00902_ ), .C1(_01323_ ), .C2(\u_reg.rf[1][26] ), .ZN(_02882_ ) );
OAI21_X1 _10039_ ( .A(_02882_ ), .B1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01341_ ), .ZN(_02883_ ) );
INV_X1 _10040_ ( .A(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02884_ ) );
OAI211_X1 _10041_ ( .A(_01327_ ), .B(_02883_ ), .C1(_02013_ ), .C2(_02884_ ), .ZN(_02885_ ) );
NAND3_X1 _10042_ ( .A1(_02881_ ), .A2(_01504_ ), .A3(_02885_ ), .ZN(_02886_ ) );
AND2_X1 _10043_ ( .A1(_02877_ ), .A2(_02886_ ), .ZN(_02887_ ) );
OAI21_X1 _10044_ ( .A(_01303_ ), .B1(_01482_ ), .B2(_02887_ ), .ZN(_02888_ ) );
AND3_X1 _10045_ ( .A1(_02292_ ), .A2(_01523_ ), .A3(_01278_ ), .ZN(_02889_ ) );
NOR3_X1 _10046_ ( .A1(_01275_ ), .A2(_01294_ ), .A3(_02889_ ), .ZN(_02890_ ) );
NAND2_X1 _10047_ ( .A1(_02890_ ), .A2(fanout_net_12 ), .ZN(_02891_ ) );
MUX2_X1 _10048_ ( .A(\ea_addr[26] ), .B(\u_exu.ecsr[26] ), .S(_01527_ ), .Z(_02892_ ) );
OR2_X1 _10049_ ( .A1(_02892_ ), .A2(fanout_net_12 ), .ZN(_02893_ ) );
AND2_X1 _10050_ ( .A1(_02891_ ), .A2(_02893_ ), .ZN(\ar_data[26] ) );
INV_X1 _10051_ ( .A(\ar_data[26] ), .ZN(_02894_ ) );
AOI21_X1 _10052_ ( .A(_02888_ ), .B1(_02894_ ), .B2(_01531_ ), .ZN(_02895_ ) );
NAND2_X1 _10053_ ( .A1(_02895_ ), .A2(_00743_ ), .ZN(_02896_ ) );
NAND4_X1 _10054_ ( .A1(_01416_ ), .A2(_00843_ ), .A3(_00842_ ), .A4(_01421_ ), .ZN(_02897_ ) );
NAND3_X1 _10055_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][26] ), .A3(_01431_ ), .ZN(_02898_ ) );
NAND3_X1 _10056_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][26] ), .A3(_01436_ ), .ZN(_02899_ ) );
NAND4_X1 _10057_ ( .A1(_02210_ ), .A2(\u_csr.csr[2][26] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_02900_ ) );
NAND3_X1 _10058_ ( .A1(_02898_ ), .A2(_02899_ ), .A3(_02900_ ), .ZN(_02901_ ) );
NAND3_X1 _10059_ ( .A1(_01537_ ), .A2(_01538_ ), .A3(_02901_ ), .ZN(_02902_ ) );
AOI21_X1 _10060_ ( .A(_01535_ ), .B1(_02897_ ), .B2(_02902_ ), .ZN(_02903_ ) );
AOI221_X4 _10061_ ( .A(_02903_ ), .B1(\de_pc[26] ), .B2(_01454_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_02904_ ) );
NAND2_X1 _10062_ ( .A1(_02895_ ), .A2(_01556_ ), .ZN(_02905_ ) );
AOI21_X1 _10063_ ( .A(_01562_ ), .B1(\u_idu.imm_auipc_lui[26] ), .B2(_01563_ ), .ZN(_02906_ ) );
NOR3_X1 _10064_ ( .A1(_02906_ ), .A2(_01555_ ), .A3(_01566_ ), .ZN(_02907_ ) );
AOI211_X1 _10065_ ( .A(_02907_ ), .B(_01052_ ), .C1(\de_pc[26] ), .C2(_01464_ ), .ZN(_02908_ ) );
AOI221_X4 _10066_ ( .A(_01644_ ), .B1(_02896_ ), .B2(_02904_ ), .C1(_02905_ ), .C2(_02908_ ), .ZN(_00156_ ) );
MUX2_X1 _10067_ ( .A(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(_01337_ ), .Z(_02909_ ) );
AND2_X1 _10068_ ( .A1(_02909_ ), .A2(_01577_ ), .ZN(_02910_ ) );
NAND3_X1 _10069_ ( .A1(_01837_ ), .A2(\u_idu.imm_auipc_lui[15] ), .A3(\u_reg.rf[1][25] ), .ZN(_02911_ ) );
AOI211_X1 _10070_ ( .A(_01484_ ), .B(_02910_ ), .C1(_01750_ ), .C2(_02911_ ), .ZN(_02912_ ) );
AOI22_X1 _10071_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01332_ ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02913_ ) );
NAND3_X1 _10072_ ( .A1(_01337_ ), .A2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01577_ ), .ZN(_02914_ ) );
NAND3_X1 _10073_ ( .A1(_01337_ ), .A2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01341_ ), .ZN(_02915_ ) );
AND4_X1 _10074_ ( .A1(_01318_ ), .A2(_02913_ ), .A3(_02914_ ), .A4(_02915_ ), .ZN(_02916_ ) );
NOR3_X1 _10075_ ( .A1(_02912_ ), .A2(_01483_ ), .A3(_02916_ ), .ZN(_02917_ ) );
AOI22_X1 _10076_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02918_ ) );
AOI22_X1 _10077_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02919_ ) );
NAND3_X1 _10078_ ( .A1(_02918_ ), .A2(_02919_ ), .A3(_01327_ ), .ZN(_02920_ ) );
AOI22_X1 _10079_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02921_ ) );
AOI22_X1 _10080_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02922_ ) );
NAND3_X1 _10081_ ( .A1(_02921_ ), .A2(_02922_ ), .A3(_01484_ ), .ZN(_02923_ ) );
AND3_X1 _10082_ ( .A1(_02920_ ), .A2(_02923_ ), .A3(_01483_ ), .ZN(_02924_ ) );
NOR2_X1 _10083_ ( .A1(_02917_ ), .A2(_02924_ ), .ZN(_02925_ ) );
OAI21_X1 _10084_ ( .A(_01303_ ), .B1(_01304_ ), .B2(_02925_ ), .ZN(_02926_ ) );
AOI21_X1 _10085_ ( .A(_01279_ ), .B1(_01887_ ), .B2(_01888_ ), .ZN(_02927_ ) );
NOR3_X1 _10086_ ( .A1(_01275_ ), .A2(_01294_ ), .A3(_02927_ ), .ZN(_02928_ ) );
NAND2_X1 _10087_ ( .A1(_02928_ ), .A2(fanout_net_12 ), .ZN(_02929_ ) );
MUX2_X1 _10088_ ( .A(\ea_addr[25] ), .B(\u_exu.ecsr[25] ), .S(_01527_ ), .Z(_02930_ ) );
OR2_X1 _10089_ ( .A1(_02930_ ), .A2(fanout_net_12 ), .ZN(_02931_ ) );
AND2_X1 _10090_ ( .A1(_02929_ ), .A2(_02931_ ), .ZN(\ar_data[25] ) );
INV_X1 _10091_ ( .A(\ar_data[25] ), .ZN(_02932_ ) );
AOI21_X1 _10092_ ( .A(_02926_ ), .B1(_02932_ ), .B2(_01531_ ), .ZN(_02933_ ) );
NAND2_X1 _10093_ ( .A1(_02933_ ), .A2(_00743_ ), .ZN(_02934_ ) );
NAND4_X1 _10094_ ( .A1(_01416_ ), .A2(_00845_ ), .A3(_00844_ ), .A4(_01421_ ), .ZN(_02935_ ) );
NAND3_X1 _10095_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][25] ), .A3(_01431_ ), .ZN(_02936_ ) );
NAND3_X1 _10096_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][25] ), .A3(_01436_ ), .ZN(_02937_ ) );
NAND4_X1 _10097_ ( .A1(_02210_ ), .A2(\u_csr.csr[2][25] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_02938_ ) );
NAND3_X1 _10098_ ( .A1(_02936_ ), .A2(_02937_ ), .A3(_02938_ ), .ZN(_02939_ ) );
NAND3_X1 _10099_ ( .A1(_01537_ ), .A2(_01538_ ), .A3(_02939_ ), .ZN(_02940_ ) );
AOI21_X1 _10100_ ( .A(_01535_ ), .B1(_02935_ ), .B2(_02940_ ), .ZN(_02941_ ) );
AOI221_X4 _10101_ ( .A(_02941_ ), .B1(\de_pc[25] ), .B2(_01454_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_02942_ ) );
NAND2_X1 _10102_ ( .A1(_02933_ ), .A2(_01556_ ), .ZN(_02943_ ) );
AOI21_X1 _10103_ ( .A(_01562_ ), .B1(\u_idu.imm_auipc_lui[25] ), .B2(_00738_ ), .ZN(_02944_ ) );
NOR3_X1 _10104_ ( .A1(_02944_ ), .A2(_01555_ ), .A3(_01565_ ), .ZN(_02945_ ) );
AOI211_X1 _10105_ ( .A(_02945_ ), .B(_01052_ ), .C1(\de_pc[25] ), .C2(_01464_ ), .ZN(_02946_ ) );
AOI221_X4 _10106_ ( .A(_00896_ ), .B1(_02934_ ), .B2(_02942_ ), .C1(_02943_ ), .C2(_02946_ ), .ZN(_00157_ ) );
AND3_X1 _10107_ ( .A1(_01959_ ), .A2(_01523_ ), .A3(_01278_ ), .ZN(_02947_ ) );
NOR3_X1 _10108_ ( .A1(_01275_ ), .A2(_01295_ ), .A3(_02947_ ), .ZN(_02948_ ) );
NAND2_X1 _10109_ ( .A1(_02948_ ), .A2(fanout_net_12 ), .ZN(_02949_ ) );
MUX2_X1 _10110_ ( .A(\ea_addr[24] ), .B(\u_exu.ecsr[24] ), .S(_01299_ ), .Z(_02950_ ) );
OR2_X1 _10111_ ( .A1(_02950_ ), .A2(fanout_net_12 ), .ZN(_02951_ ) );
AOI21_X1 _10112_ ( .A(_01245_ ), .B1(_02949_ ), .B2(_02951_ ), .ZN(_02952_ ) );
AOI22_X1 _10113_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02953_ ) );
AOI22_X1 _10114_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02954_ ) );
NAND3_X1 _10115_ ( .A1(_02953_ ), .A2(_02954_ ), .A3(_01312_ ), .ZN(_02955_ ) );
AOI22_X1 _10116_ ( .A1(_01005_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01314_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02956_ ) );
AOI22_X1 _10117_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01306_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02957_ ) );
NAND3_X1 _10118_ ( .A1(_02956_ ), .A2(_02957_ ), .A3(_00915_ ), .ZN(_02958_ ) );
AND3_X1 _10119_ ( .A1(_02955_ ), .A2(_02958_ ), .A3(_01320_ ), .ZN(_02959_ ) );
NAND3_X1 _10120_ ( .A1(_01338_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01339_ ), .ZN(_02960_ ) );
INV_X1 _10121_ ( .A(\u_reg.rf[1][24] ), .ZN(_02961_ ) );
AOI21_X1 _10122_ ( .A(_01506_ ), .B1(_01342_ ), .B2(_02961_ ), .ZN(_02962_ ) );
NOR2_X1 _10123_ ( .A1(_01589_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02963_ ) );
OAI211_X1 _10124_ ( .A(_01580_ ), .B(_02960_ ), .C1(_02962_ ), .C2(_02963_ ), .ZN(_02964_ ) );
AOI22_X1 _10125_ ( .A1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01495_ ), .B1(_01492_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02965_ ) );
NAND3_X1 _10126_ ( .A1(_01337_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01577_ ), .ZN(_02966_ ) );
NAND3_X1 _10127_ ( .A1(_01337_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01341_ ), .ZN(_02967_ ) );
NAND4_X1 _10128_ ( .A1(_02965_ ), .A2(_01318_ ), .A3(_02966_ ), .A4(_02967_ ), .ZN(_02968_ ) );
AND2_X1 _10129_ ( .A1(_02968_ ), .A2(_01046_ ), .ZN(_02969_ ) );
AOI21_X1 _10130_ ( .A(_02959_ ), .B1(_02964_ ), .B2(_02969_ ), .ZN(_02970_ ) );
OAI21_X1 _10131_ ( .A(_00736_ ), .B1(_01304_ ), .B2(_02970_ ), .ZN(_02971_ ) );
OR3_X1 _10132_ ( .A1(_02952_ ), .A2(_00723_ ), .A3(_02971_ ), .ZN(_02972_ ) );
AND4_X1 _10133_ ( .A1(\u_csr.csr[2][24] ), .A2(_01539_ ), .A3(_01620_ ), .A4(_01622_ ), .ZN(_02973_ ) );
NOR3_X1 _10134_ ( .A1(_02973_ ), .A2(_01544_ ), .A3(_01627_ ), .ZN(_02974_ ) );
AND4_X1 _10135_ ( .A1(\u_csr.csr[0][24] ), .A2(_01439_ ), .A3(_01410_ ), .A4(_01548_ ), .ZN(_02975_ ) );
AOI21_X1 _10136_ ( .A(_02975_ ), .B1(_01631_ ), .B2(\u_csr.csr[1][24] ), .ZN(_02976_ ) );
AOI21_X1 _10137_ ( .A(_01619_ ), .B1(_02974_ ), .B2(_02976_ ), .ZN(_02977_ ) );
AOI211_X1 _10138_ ( .A(_01419_ ), .B(_01537_ ), .C1(_00846_ ), .C2(_00847_ ), .ZN(_02978_ ) );
NOR2_X1 _10139_ ( .A1(_02977_ ), .A2(_02978_ ), .ZN(_02979_ ) );
NOR2_X1 _10140_ ( .A1(_02979_ ), .A2(_01353_ ), .ZN(_02980_ ) );
AOI211_X1 _10141_ ( .A(_01050_ ), .B(_02980_ ), .C1(\de_pc[24] ), .C2(_01455_ ), .ZN(_02981_ ) );
OR3_X1 _10142_ ( .A1(_02952_ ), .A2(_01460_ ), .A3(_02971_ ), .ZN(_02982_ ) );
AOI21_X1 _10143_ ( .A(_01562_ ), .B1(\u_idu.imm_auipc_lui[24] ), .B2(_00738_ ), .ZN(_02983_ ) );
NOR3_X1 _10144_ ( .A1(_02983_ ), .A2(_01555_ ), .A3(_01565_ ), .ZN(_02984_ ) );
AOI211_X1 _10145_ ( .A(_02984_ ), .B(_01052_ ), .C1(\de_pc[24] ), .C2(_01464_ ), .ZN(_02985_ ) );
AOI221_X1 _10146_ ( .A(_00896_ ), .B1(_02972_ ), .B2(_02981_ ), .C1(_02982_ ), .C2(_02985_ ), .ZN(_00158_ ) );
AOI22_X1 _10147_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02986_ ) );
AOI22_X1 _10148_ ( .A1(_01570_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02987_ ) );
NAND3_X1 _10149_ ( .A1(_02986_ ), .A2(_02987_ ), .A3(_01312_ ), .ZN(_02988_ ) );
AOI22_X1 _10150_ ( .A1(_01308_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01310_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02989_ ) );
AOI22_X1 _10151_ ( .A1(_01305_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01332_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02990_ ) );
NAND3_X1 _10152_ ( .A1(_02989_ ), .A2(_02990_ ), .A3(_01318_ ), .ZN(_02991_ ) );
AND3_X1 _10153_ ( .A1(_02988_ ), .A2(_02991_ ), .A3(_01320_ ), .ZN(_02992_ ) );
NAND3_X1 _10154_ ( .A1(_01586_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01587_ ), .ZN(_02993_ ) );
INV_X1 _10155_ ( .A(\u_reg.rf[1][23] ), .ZN(_02994_ ) );
AOI21_X1 _10156_ ( .A(_01506_ ), .B1(_01589_ ), .B2(_02994_ ), .ZN(_02995_ ) );
NOR2_X1 _10157_ ( .A1(_01589_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02996_ ) );
OAI211_X1 _10158_ ( .A(_01580_ ), .B(_02993_ ), .C1(_02995_ ), .C2(_02996_ ), .ZN(_02997_ ) );
AOI22_X1 _10159_ ( .A1(_01494_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01495_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02998_ ) );
AOI22_X1 _10160_ ( .A1(_01488_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02999_ ) );
NAND3_X1 _10161_ ( .A1(_02998_ ), .A2(_02999_ ), .A3(_01336_ ), .ZN(_03000_ ) );
AND2_X1 _10162_ ( .A1(_03000_ ), .A2(_01046_ ), .ZN(_03001_ ) );
AOI21_X1 _10163_ ( .A(_02992_ ), .B1(_02997_ ), .B2(_03001_ ), .ZN(_03002_ ) );
OAI21_X1 _10164_ ( .A(_01303_ ), .B1(_01304_ ), .B2(_03002_ ), .ZN(_03003_ ) );
AOI21_X1 _10165_ ( .A(_01884_ ), .B1(_01261_ ), .B2(_01262_ ), .ZN(_03004_ ) );
MUX2_X1 _10166_ ( .A(_03004_ ), .B(_01269_ ), .S(_01523_ ), .Z(_03005_ ) );
AOI21_X1 _10167_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_03005_ ), .ZN(_03006_ ) );
NAND2_X1 _10168_ ( .A1(_03006_ ), .A2(fanout_net_12 ), .ZN(_03007_ ) );
MUX2_X1 _10169_ ( .A(\ea_addr[23] ), .B(\u_exu.ecsr[23] ), .S(_01527_ ), .Z(_03008_ ) );
OR2_X1 _10170_ ( .A1(_03008_ ), .A2(\u_arbiter.rvalid ), .ZN(_03009_ ) );
AND2_X1 _10171_ ( .A1(_03007_ ), .A2(_03009_ ), .ZN(\ar_data[23] ) );
INV_X1 _10172_ ( .A(\ar_data[23] ), .ZN(_03010_ ) );
AOI21_X2 _10173_ ( .A(_03003_ ), .B1(_03010_ ), .B2(_01482_ ), .ZN(_03011_ ) );
NAND2_X1 _10174_ ( .A1(_03011_ ), .A2(_00743_ ), .ZN(_03012_ ) );
NAND4_X1 _10175_ ( .A1(_01416_ ), .A2(_00849_ ), .A3(_00848_ ), .A4(_01421_ ), .ZN(_03013_ ) );
NAND3_X1 _10176_ ( .A1(_01429_ ), .A2(\u_csr.csr[1][23] ), .A3(_01431_ ), .ZN(_03014_ ) );
NAND3_X1 _10177_ ( .A1(_01434_ ), .A2(\u_csr.csr[0][23] ), .A3(_01436_ ), .ZN(_03015_ ) );
NAND4_X1 _10178_ ( .A1(_02210_ ), .A2(\u_csr.csr[2][23] ), .A3(_01440_ ), .A4(_01442_ ), .ZN(_03016_ ) );
NAND3_X1 _10179_ ( .A1(_03014_ ), .A2(_03015_ ), .A3(_03016_ ), .ZN(_03017_ ) );
NAND3_X1 _10180_ ( .A1(_01537_ ), .A2(_01538_ ), .A3(_03017_ ), .ZN(_03018_ ) );
AOI21_X1 _10181_ ( .A(_01352_ ), .B1(_03013_ ), .B2(_03018_ ), .ZN(_03019_ ) );
AOI221_X4 _10182_ ( .A(_03019_ ), .B1(\de_pc[23] ), .B2(_01454_ ), .C1(_01062_ ), .C2(_01065_ ), .ZN(_03020_ ) );
NAND2_X1 _10183_ ( .A1(_03011_ ), .A2(_01556_ ), .ZN(_03021_ ) );
OAI21_X1 _10184_ ( .A(_01561_ ), .B1(_00893_ ), .B2(_00928_ ), .ZN(_03022_ ) );
AOI221_X4 _10185_ ( .A(_01051_ ), .B1(\de_pc[23] ), .B2(_01463_ ), .C1(_01467_ ), .C2(_03022_ ), .ZN(_03023_ ) );
AOI221_X1 _10186_ ( .A(_00896_ ), .B1(_03012_ ), .B2(_03020_ ), .C1(_03021_ ), .C2(_03023_ ), .ZN(_00159_ ) );
AOI22_X1 _10187_ ( .A1(_01316_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_00909_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03024_ ) );
AOI22_X1 _10188_ ( .A1(_01005_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01309_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03025_ ) );
NAND3_X1 _10189_ ( .A1(_03024_ ), .A2(_03025_ ), .A3(_00975_ ), .ZN(_03026_ ) );
AOI22_X1 _10190_ ( .A1(_01005_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01309_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03027_ ) );
AOI22_X1 _10191_ ( .A1(_00950_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_00909_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03028_ ) );
NAND3_X1 _10192_ ( .A1(_03027_ ), .A2(_03028_ ), .A3(_00915_ ), .ZN(_03029_ ) );
AND3_X1 _10193_ ( .A1(_03026_ ), .A2(_03029_ ), .A3(_01320_ ), .ZN(_03030_ ) );
OAI211_X1 _10194_ ( .A(\u_idu.imm_auipc_lui[15] ), .B(_00902_ ), .C1(_01323_ ), .C2(\u_reg.rf[1][22] ), .ZN(_03031_ ) );
OAI21_X1 _10195_ ( .A(_03031_ ), .B1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01341_ ), .ZN(_03032_ ) );
NAND4_X1 _10196_ ( .A1(_01323_ ), .A2(\u_idu.imm_auipc_lui[15] ), .A3(_00902_ ), .A4(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03033_ ) );
NAND3_X1 _10197_ ( .A1(_03032_ ), .A2(_00975_ ), .A3(_03033_ ), .ZN(_03034_ ) );
AND2_X1 _10198_ ( .A1(_03034_ ), .A2(_01046_ ), .ZN(_03035_ ) );
AOI22_X1 _10199_ ( .A1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01486_ ), .B1(_01489_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03036_ ) );
NAND3_X1 _10200_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01328_ ), .ZN(_03037_ ) );
NAND3_X1 _10201_ ( .A1(_01500_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01325_ ), .ZN(_03038_ ) );
NAND4_X1 _10202_ ( .A1(_03036_ ), .A2(_01484_ ), .A3(_03037_ ), .A4(_03038_ ), .ZN(_03039_ ) );
AOI21_X1 _10203_ ( .A(_03030_ ), .B1(_03035_ ), .B2(_03039_ ), .ZN(_03040_ ) );
OAI21_X1 _10204_ ( .A(_00736_ ), .B1(_01244_ ), .B2(_03040_ ), .ZN(_03041_ ) );
AND3_X1 _10205_ ( .A1(_01514_ ), .A2(_01270_ ), .A3(_01521_ ), .ZN(_03042_ ) );
MUX2_X1 _10206_ ( .A(_02067_ ), .B(_03042_ ), .S(_01253_ ), .Z(_03043_ ) );
AOI21_X1 _10207_ ( .A(_01594_ ), .B1(\io_master_arsize[1] ), .B2(_03043_ ), .ZN(_03044_ ) );
NAND2_X1 _10208_ ( .A1(_03044_ ), .A2(\u_arbiter.rvalid ), .ZN(_03045_ ) );
MUX2_X1 _10209_ ( .A(\ea_addr[22] ), .B(\u_exu.ecsr[22] ), .S(_01298_ ), .Z(_03046_ ) );
OR2_X1 _10210_ ( .A1(_03046_ ), .A2(\u_arbiter.rvalid ), .ZN(_03047_ ) );
AND2_X1 _10211_ ( .A1(_03045_ ), .A2(_03047_ ), .ZN(\ar_data[22] ) );
INV_X1 _10212_ ( .A(\ar_data[22] ), .ZN(_03048_ ) );
AOI21_X1 _10213_ ( .A(_03041_ ), .B1(_03048_ ), .B2(_01304_ ), .ZN(_03049_ ) );
NAND2_X1 _10214_ ( .A1(_03049_ ), .A2(_01556_ ), .ZN(_03050_ ) );
OAI21_X1 _10215_ ( .A(_01561_ ), .B1(_00894_ ), .B2(_00928_ ), .ZN(_03051_ ) );
AOI221_X4 _10216_ ( .A(_01051_ ), .B1(\de_pc[22] ), .B2(_01463_ ), .C1(_01467_ ), .C2(_03051_ ), .ZN(_03052_ ) );
NAND2_X1 _10217_ ( .A1(_03049_ ), .A2(_00743_ ), .ZN(_03053_ ) );
INV_X1 _10218_ ( .A(_01450_ ), .ZN(_03054_ ) );
NAND3_X1 _10219_ ( .A1(_03054_ ), .A2(\de_pc[22] ), .A3(_00723_ ), .ZN(_03055_ ) );
NAND2_X1 _10220_ ( .A1(_03053_ ), .A2(_03055_ ), .ZN(_03056_ ) );
AND3_X1 _10221_ ( .A1(_01433_ ), .A2(\u_csr.csr[0][22] ), .A3(_01435_ ), .ZN(_03057_ ) );
NAND4_X1 _10222_ ( .A1(_01539_ ), .A2(\u_csr.csr[2][22] ), .A3(_00755_ ), .A4(_01621_ ), .ZN(_03058_ ) );
NAND3_X1 _10223_ ( .A1(_01545_ ), .A2(_01692_ ), .A3(_03058_ ), .ZN(_03059_ ) );
AOI211_X1 _10224_ ( .A(_03057_ ), .B(_03059_ ), .C1(\u_csr.csr[1][22] ), .C2(_01631_ ), .ZN(_03060_ ) );
OR2_X1 _10225_ ( .A1(_01619_ ), .A2(_03060_ ), .ZN(_03061_ ) );
NAND4_X1 _10226_ ( .A1(_01713_ ), .A2(_00851_ ), .A3(_00850_ ), .A4(_01425_ ), .ZN(_03062_ ) );
AND2_X1 _10227_ ( .A1(_03061_ ), .A2(_03062_ ), .ZN(_03063_ ) );
OR2_X1 _10228_ ( .A1(_03063_ ), .A2(_00758_ ), .ZN(_03064_ ) );
INV_X1 _10229_ ( .A(\de_pc[22] ), .ZN(_03065_ ) );
INV_X1 _10230_ ( .A(_00758_ ), .ZN(_03066_ ) );
OAI21_X1 _10231_ ( .A(_03064_ ), .B1(_03065_ ), .B2(_03066_ ), .ZN(_03067_ ) );
AOI21_X1 _10232_ ( .A(_03056_ ), .B1(_01450_ ), .B2(_03067_ ), .ZN(_03068_ ) );
AOI221_X1 _10233_ ( .A(_00896_ ), .B1(_03050_ ), .B2(_03052_ ), .C1(_03068_ ), .C2(_01053_ ), .ZN(_00160_ ) );
NOR2_X1 _10234_ ( .A1(\u_exu.alu_ctrl[5] ), .A2(\u_exu.alu_ctrl[4] ), .ZN(_03069_ ) );
AND2_X2 _10235_ ( .A1(_03069_ ), .A2(fanout_net_20 ), .ZN(_03070_ ) );
INV_X2 _10236_ ( .A(_03070_ ), .ZN(_03071_ ) );
INV_X32 _10237_ ( .A(\u_exu.alu_ctrl[3] ), .ZN(_03072_ ) );
BUF_X32 _10238_ ( .A(_03072_ ), .Z(_03073_ ) );
BUF_X4 _10239_ ( .A(_03073_ ), .Z(_03074_ ) );
BUF_X16 _10240_ ( .A(_03074_ ), .Z(_03075_ ) );
AND3_X1 _10241_ ( .A1(_03075_ ), .A2(fanout_net_13 ), .A3(\u_exu.alu_p1[0] ), .ZN(_03076_ ) );
INV_X1 _10242_ ( .A(\u_exu.alu_ctrl[4] ), .ZN(_03077_ ) );
NOR2_X1 _10243_ ( .A1(_03077_ ), .A2(\u_exu.alu_ctrl[5] ), .ZN(_03078_ ) );
INV_X1 _10244_ ( .A(fanout_net_13 ), .ZN(_03079_ ) );
CLKBUF_X2 _10245_ ( .A(_03079_ ), .Z(_03080_ ) );
NOR2_X1 _10246_ ( .A1(_03080_ ), .A2(\u_exu.alu_ctrl[3] ), .ZN(_03081_ ) );
OAI211_X1 _10247_ ( .A(fanout_net_20 ), .B(_03078_ ), .C1(_03081_ ), .C2(\u_exu.alu_p1[0] ), .ZN(_03082_ ) );
AND2_X1 _10248_ ( .A1(\u_exu.alu_ctrl[5] ), .A2(\u_exu.alu_ctrl[4] ), .ZN(_03083_ ) );
AND2_X1 _10249_ ( .A1(_03083_ ), .A2(fanout_net_20 ), .ZN(_03084_ ) );
XOR2_X1 _10250_ ( .A(\u_exu.alu_p2[4] ), .B(\u_exu.alu_p1[4] ), .Z(_03085_ ) );
XOR2_X1 _10251_ ( .A(fanout_net_15 ), .B(\u_exu.alu_p1[1] ), .Z(_03086_ ) );
XOR2_X1 _10252_ ( .A(\u_exu.alu_p1[7] ), .B(\u_exu.alu_p2[7] ), .Z(_03087_ ) );
AND2_X1 _10253_ ( .A1(fanout_net_17 ), .A2(\u_exu.alu_p1[2] ), .ZN(_03088_ ) );
NOR2_X1 _10254_ ( .A1(fanout_net_17 ), .A2(\u_exu.alu_p1[2] ), .ZN(_03089_ ) );
NOR2_X1 _10255_ ( .A1(_03088_ ), .A2(_03089_ ), .ZN(_03090_ ) );
NOR4_X1 _10256_ ( .A1(_03085_ ), .A2(_03086_ ), .A3(_03087_ ), .A4(_03090_ ), .ZN(_03091_ ) );
XOR2_X1 _10257_ ( .A(\u_exu.alu_p1[12] ), .B(\u_exu.alu_p2[12] ), .Z(_03092_ ) );
XOR2_X1 _10258_ ( .A(\u_exu.alu_p1[10] ), .B(\u_exu.alu_p2[10] ), .Z(_03093_ ) );
XOR2_X1 _10259_ ( .A(\u_exu.alu_p2[9] ), .B(\u_exu.alu_p1[9] ), .Z(_03094_ ) );
XOR2_X1 _10260_ ( .A(\u_exu.alu_p1[15] ), .B(\u_exu.alu_p2[15] ), .Z(_03095_ ) );
NOR4_X1 _10261_ ( .A1(_03092_ ), .A2(_03093_ ), .A3(_03094_ ), .A4(_03095_ ), .ZN(_03096_ ) );
XOR2_X1 _10262_ ( .A(\u_exu.alu_p1[26] ), .B(\u_exu.alu_p2[26] ), .Z(_03097_ ) );
XOR2_X1 _10263_ ( .A(\u_exu.alu_p1[31] ), .B(\u_exu.alu_p2[31] ), .Z(_03098_ ) );
XOR2_X1 _10264_ ( .A(\u_exu.alu_p1[28] ), .B(\u_exu.alu_p2[28] ), .Z(_03099_ ) );
XOR2_X1 _10265_ ( .A(\u_exu.alu_p1[25] ), .B(\u_exu.alu_p2[25] ), .Z(_03100_ ) );
NOR4_X1 _10266_ ( .A1(_03097_ ), .A2(_03098_ ), .A3(_03099_ ), .A4(_03100_ ), .ZN(_03101_ ) );
XOR2_X1 _10267_ ( .A(\u_exu.alu_p1[20] ), .B(\u_exu.alu_p2[20] ), .Z(_03102_ ) );
XOR2_X1 _10268_ ( .A(\u_exu.alu_p1[19] ), .B(\u_exu.alu_p2[19] ), .Z(_03103_ ) );
XOR2_X1 _10269_ ( .A(\u_exu.alu_p1[22] ), .B(\u_exu.alu_p2[22] ), .Z(_03104_ ) );
AND2_X1 _10270_ ( .A1(\u_exu.alu_p1[16] ), .A2(\u_exu.alu_p2[16] ), .ZN(_03105_ ) );
NOR2_X1 _10271_ ( .A1(\u_exu.alu_p1[16] ), .A2(\u_exu.alu_p2[16] ), .ZN(_03106_ ) );
NOR2_X1 _10272_ ( .A1(_03105_ ), .A2(_03106_ ), .ZN(_03107_ ) );
NOR4_X1 _10273_ ( .A1(_03102_ ), .A2(_03103_ ), .A3(_03104_ ), .A4(_03107_ ), .ZN(_03108_ ) );
AND4_X1 _10274_ ( .A1(_03091_ ), .A2(_03096_ ), .A3(_03101_ ), .A4(_03108_ ), .ZN(_03109_ ) );
XOR2_X1 _10275_ ( .A(fanout_net_13 ), .B(\u_exu.alu_p1[0] ), .Z(_03110_ ) );
XOR2_X1 _10276_ ( .A(\u_exu.alu_p1[6] ), .B(\u_exu.alu_p2[6] ), .Z(_03111_ ) );
XOR2_X1 _10277_ ( .A(fanout_net_19 ), .B(\u_exu.alu_p1[3] ), .Z(_03112_ ) );
XOR2_X1 _10278_ ( .A(\u_exu.alu_p1[5] ), .B(\u_exu.alu_p2[5] ), .Z(_03113_ ) );
NOR4_X1 _10279_ ( .A1(_03110_ ), .A2(_03111_ ), .A3(_03112_ ), .A4(_03113_ ), .ZN(_03114_ ) );
XOR2_X1 _10280_ ( .A(\u_exu.alu_p1[13] ), .B(\u_exu.alu_p2[13] ), .Z(_03115_ ) );
XOR2_X1 _10281_ ( .A(\u_exu.alu_p1[8] ), .B(\u_exu.alu_p2[8] ), .Z(_03116_ ) );
XOR2_X1 _10282_ ( .A(\u_exu.alu_p1[14] ), .B(\u_exu.alu_p2[14] ), .Z(_03117_ ) );
XOR2_X1 _10283_ ( .A(\u_exu.alu_p1[11] ), .B(\u_exu.alu_p2[11] ), .Z(_03118_ ) );
NOR4_X1 _10284_ ( .A1(_03115_ ), .A2(_03116_ ), .A3(_03117_ ), .A4(_03118_ ), .ZN(_03119_ ) );
XOR2_X1 _10285_ ( .A(\u_exu.alu_p2[17] ), .B(\u_exu.alu_p1[17] ), .Z(_03120_ ) );
XOR2_X1 _10286_ ( .A(\u_exu.alu_p1[18] ), .B(\u_exu.alu_p2[18] ), .Z(_03121_ ) );
XOR2_X1 _10287_ ( .A(\u_exu.alu_p1[21] ), .B(\u_exu.alu_p2[21] ), .Z(_03122_ ) );
XOR2_X1 _10288_ ( .A(\u_exu.alu_p1[23] ), .B(\u_exu.alu_p2[23] ), .Z(_03123_ ) );
NOR4_X1 _10289_ ( .A1(_03120_ ), .A2(_03121_ ), .A3(_03122_ ), .A4(_03123_ ), .ZN(_03124_ ) );
XOR2_X1 _10290_ ( .A(\u_exu.alu_p1[30] ), .B(\u_exu.alu_p2[30] ), .Z(_03125_ ) );
XOR2_X1 _10291_ ( .A(\u_exu.alu_p1[27] ), .B(\u_exu.alu_p2[27] ), .Z(_03126_ ) );
XOR2_X1 _10292_ ( .A(\u_exu.alu_p1[24] ), .B(\u_exu.alu_p2[24] ), .Z(_03127_ ) );
AND2_X1 _10293_ ( .A1(\u_exu.alu_p1[29] ), .A2(\u_exu.alu_p2[29] ), .ZN(_03128_ ) );
NOR2_X1 _10294_ ( .A1(\u_exu.alu_p1[29] ), .A2(\u_exu.alu_p2[29] ), .ZN(_03129_ ) );
NOR2_X1 _10295_ ( .A1(_03128_ ), .A2(_03129_ ), .ZN(_03130_ ) );
NOR4_X1 _10296_ ( .A1(_03125_ ), .A2(_03126_ ), .A3(_03127_ ), .A4(_03130_ ), .ZN(_03131_ ) );
AND4_X1 _10297_ ( .A1(_03114_ ), .A2(_03119_ ), .A3(_03124_ ), .A4(_03131_ ), .ZN(_03132_ ) );
NAND3_X1 _10298_ ( .A1(_03109_ ), .A2(_03132_ ), .A3(\u_exu.alu_ctrl[2] ), .ZN(_03133_ ) );
AND3_X1 _10299_ ( .A1(\u_exu.alu_ctrl[6] ), .A2(\u_exu.alu_ctrl[5] ), .A3(\u_exu.alu_ctrl[4] ), .ZN(_03134_ ) );
AND2_X1 _10300_ ( .A1(_03133_ ), .A2(_03134_ ), .ZN(_03135_ ) );
AND2_X1 _10301_ ( .A1(_03109_ ), .A2(_03132_ ), .ZN(_03136_ ) );
OAI21_X1 _10302_ ( .A(_03135_ ), .B1(\u_exu.alu_ctrl[2] ), .B2(_03136_ ), .ZN(_03137_ ) );
NAND2_X1 _10303_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[30] ), .ZN(_03138_ ) );
INV_X32 _10304_ ( .A(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03139_ ) );
BUF_X32 _10305_ ( .A(_03139_ ), .Z(_03140_ ) );
BUF_X32 _10306_ ( .A(_03140_ ), .Z(_03141_ ) );
BUF_X4 _10307_ ( .A(_03141_ ), .Z(_03142_ ) );
XNOR2_X1 _10308_ ( .A(_03138_ ), .B(_03142_ ), .ZN(_03143_ ) );
INV_X1 _10309_ ( .A(\u_exu.alu_p1[30] ), .ZN(_03144_ ) );
XNOR2_X1 _10310_ ( .A(_03143_ ), .B(_03144_ ), .ZN(_03145_ ) );
INV_X1 _10311_ ( .A(_03145_ ), .ZN(_03146_ ) );
NAND2_X4 _10312_ ( .A1(_03073_ ), .A2(\u_exu.alu_p2[15] ), .ZN(_03147_ ) );
XNOR2_X2 _10313_ ( .A(_03147_ ), .B(_03140_ ), .ZN(_03148_ ) );
XNOR2_X2 _10314_ ( .A(_03148_ ), .B(\u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03149_ ) );
NAND2_X1 _10315_ ( .A1(_03073_ ), .A2(\u_exu.alu_p2[14] ), .ZN(_03150_ ) );
XNOR2_X2 _10316_ ( .A(_03150_ ), .B(_03141_ ), .ZN(_03151_ ) );
AND2_X1 _10317_ ( .A1(_03151_ ), .A2(\u_exu.alu_p1[14] ), .ZN(_03152_ ) );
AND2_X1 _10318_ ( .A1(_03149_ ), .A2(_03152_ ), .ZN(_03153_ ) );
NAND2_X1 _10319_ ( .A1(_03072_ ), .A2(\u_exu.alu_p2[11] ), .ZN(_03154_ ) );
NAND2_X1 _10320_ ( .A1(_03154_ ), .A2(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03155_ ) );
NAND3_X4 _10321_ ( .A1(_03140_ ), .A2(_03073_ ), .A3(\u_exu.alu_p2[11] ), .ZN(_03156_ ) );
AND2_X4 _10322_ ( .A1(_03155_ ), .A2(_03156_ ), .ZN(_03157_ ) );
XNOR2_X2 _10323_ ( .A(_03157_ ), .B(\u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03158_ ) );
NAND2_X4 _10324_ ( .A1(_03073_ ), .A2(\u_exu.alu_p2[10] ), .ZN(_03159_ ) );
XNOR2_X2 _10325_ ( .A(_03159_ ), .B(_03140_ ), .ZN(_03160_ ) );
AND2_X1 _10326_ ( .A1(_03160_ ), .A2(\u_exu.alu_p1[10] ), .ZN(_03161_ ) );
NAND2_X1 _10327_ ( .A1(_03158_ ), .A2(_03161_ ), .ZN(_03162_ ) );
INV_X1 _10328_ ( .A(_03157_ ), .ZN(_03163_ ) );
OAI21_X1 _10329_ ( .A(_03162_ ), .B1(\u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B2(_03163_ ), .ZN(_03164_ ) );
NAND2_X4 _10330_ ( .A1(_03072_ ), .A2(\u_exu.alu_p2[9] ), .ZN(_03165_ ) );
XNOR2_X2 _10331_ ( .A(_03165_ ), .B(_03139_ ), .ZN(_03166_ ) );
XNOR2_X2 _10332_ ( .A(_03166_ ), .B(\u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03167_ ) );
NAND2_X4 _10333_ ( .A1(_03072_ ), .A2(\u_exu.alu_p2[8] ), .ZN(_03168_ ) );
XNOR2_X1 _10334_ ( .A(_03168_ ), .B(_03139_ ), .ZN(_03169_ ) );
AND2_X4 _10335_ ( .A1(_03169_ ), .A2(\u_exu.alu_p1[8] ), .ZN(_03170_ ) );
AND2_X4 _10336_ ( .A1(_03167_ ), .A2(_03170_ ), .ZN(_03171_ ) );
INV_X1 _10337_ ( .A(\u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03172_ ) );
AOI21_X2 _10338_ ( .A(_03171_ ), .B1(_03172_ ), .B2(_03166_ ), .ZN(_03173_ ) );
INV_X2 _10339_ ( .A(_03173_ ), .ZN(_03174_ ) );
INV_X1 _10340_ ( .A(\u_exu.alu_p1[10] ), .ZN(_03175_ ) );
XNOR2_X2 _10341_ ( .A(_03160_ ), .B(_03175_ ), .ZN(_03176_ ) );
AND2_X2 _10342_ ( .A1(_03176_ ), .A2(_03158_ ), .ZN(_03177_ ) );
AOI21_X4 _10343_ ( .A(_03164_ ), .B1(_03174_ ), .B2(_03177_ ), .ZN(_03178_ ) );
INV_X1 _10344_ ( .A(\u_exu.alu_p1[14] ), .ZN(_03179_ ) );
XNOR2_X2 _10345_ ( .A(_03151_ ), .B(_03179_ ), .ZN(_03180_ ) );
AND2_X2 _10346_ ( .A1(_03180_ ), .A2(_03149_ ), .ZN(_03181_ ) );
NAND2_X4 _10347_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[12] ), .ZN(_03182_ ) );
XNOR2_X2 _10348_ ( .A(_03182_ ), .B(_03141_ ), .ZN(_03183_ ) );
INV_X1 _10349_ ( .A(\u_exu.alu_p1[12] ), .ZN(_03184_ ) );
XNOR2_X1 _10350_ ( .A(_03183_ ), .B(_03184_ ), .ZN(_03185_ ) );
NAND2_X4 _10351_ ( .A1(_03073_ ), .A2(\u_exu.alu_p2[13] ), .ZN(_03186_ ) );
XNOR2_X1 _10352_ ( .A(_03186_ ), .B(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03187_ ) );
XNOR2_X2 _10353_ ( .A(_03187_ ), .B(\u_exu.alu_p1[13] ), .ZN(_03188_ ) );
NAND3_X2 _10354_ ( .A1(_03181_ ), .A2(_03185_ ), .A3(_03188_ ), .ZN(_03189_ ) );
NOR2_X2 _10355_ ( .A1(_03178_ ), .A2(_03189_ ), .ZN(_03190_ ) );
INV_X1 _10356_ ( .A(_03181_ ), .ZN(_03191_ ) );
INV_X1 _10357_ ( .A(\u_exu.alu_p1[13] ), .ZN(_03192_ ) );
NOR2_X1 _10358_ ( .A1(_03187_ ), .A2(_03192_ ), .ZN(_03193_ ) );
INV_X1 _10359_ ( .A(_03193_ ), .ZN(_03194_ ) );
AND2_X1 _10360_ ( .A1(_03183_ ), .A2(\u_exu.alu_p1[12] ), .ZN(_03195_ ) );
NAND2_X1 _10361_ ( .A1(_03188_ ), .A2(_03195_ ), .ZN(_03196_ ) );
AOI21_X2 _10362_ ( .A(_03191_ ), .B1(_03194_ ), .B2(_03196_ ), .ZN(_03197_ ) );
OR2_X4 _10363_ ( .A1(_03190_ ), .A2(_03197_ ), .ZN(_03198_ ) );
INV_X1 _10364_ ( .A(\u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03199_ ) );
AOI211_X2 _10365_ ( .A(_03153_ ), .B(_03198_ ), .C1(_03199_ ), .C2(_03148_ ), .ZN(_03200_ ) );
NAND2_X4 _10366_ ( .A1(_03073_ ), .A2(\u_exu.alu_p2[6] ), .ZN(_03201_ ) );
XNOR2_X2 _10367_ ( .A(_03201_ ), .B(_03140_ ), .ZN(_03202_ ) );
INV_X1 _10368_ ( .A(\u_exu.alu_p1[6] ), .ZN(_03203_ ) );
XNOR2_X2 _10369_ ( .A(_03202_ ), .B(_03203_ ), .ZN(_03204_ ) );
NAND2_X4 _10370_ ( .A1(_03073_ ), .A2(\u_exu.alu_p2[7] ), .ZN(_03205_ ) );
NAND2_X4 _10371_ ( .A1(_03205_ ), .A2(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03206_ ) );
NAND3_X4 _10372_ ( .A1(_03140_ ), .A2(_03073_ ), .A3(\u_exu.alu_p2[7] ), .ZN(_03207_ ) );
AND2_X4 _10373_ ( .A1(_03206_ ), .A2(_03207_ ), .ZN(_03208_ ) );
XNOR2_X2 _10374_ ( .A(_03208_ ), .B(\u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03209_ ) );
NAND2_X4 _10375_ ( .A1(_03204_ ), .A2(_03209_ ), .ZN(_03210_ ) );
NAND2_X4 _10376_ ( .A1(_03073_ ), .A2(\u_exu.alu_p2[4] ), .ZN(_03211_ ) );
XNOR2_X2 _10377_ ( .A(_03211_ ), .B(_03140_ ), .ZN(_03212_ ) );
INV_X1 _10378_ ( .A(\u_exu.alu_p1[4] ), .ZN(_03213_ ) );
XNOR2_X2 _10379_ ( .A(_03212_ ), .B(_03213_ ), .ZN(_03214_ ) );
NAND2_X1 _10380_ ( .A1(_03072_ ), .A2(\u_exu.alu_p2[5] ), .ZN(_03215_ ) );
XNOR2_X2 _10381_ ( .A(_03215_ ), .B(_03140_ ), .ZN(_03216_ ) );
XNOR2_X2 _10382_ ( .A(_03216_ ), .B(\u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03217_ ) );
AND2_X4 _10383_ ( .A1(_03214_ ), .A2(_03217_ ), .ZN(_03218_ ) );
INV_X2 _10384_ ( .A(_03218_ ), .ZN(_03219_ ) );
NAND2_X1 _10385_ ( .A1(_03072_ ), .A2(fanout_net_19 ), .ZN(_03220_ ) );
XNOR2_X2 _10386_ ( .A(_03220_ ), .B(_03140_ ), .ZN(_03221_ ) );
XNOR2_X2 _10387_ ( .A(_03221_ ), .B(\u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03222_ ) );
NOR2_X4 _10388_ ( .A1(\u_exu.alu_ctrl[3] ), .A2(fanout_net_17 ), .ZN(_03223_ ) );
XNOR2_X1 _10389_ ( .A(_03223_ ), .B(\u_exu.alu_ctrl[0] ), .ZN(_03224_ ) );
INV_X1 _10390_ ( .A(\u_exu.alu_p1[2] ), .ZN(_03225_ ) );
XNOR2_X1 _10391_ ( .A(_03224_ ), .B(_03225_ ), .ZN(_03226_ ) );
NAND2_X1 _10392_ ( .A1(_03072_ ), .A2(fanout_net_15 ), .ZN(_03227_ ) );
XNOR2_X2 _10393_ ( .A(_03227_ ), .B(_03140_ ), .ZN(_03228_ ) );
XNOR2_X2 _10394_ ( .A(_03228_ ), .B(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ), .ZN(_03229_ ) );
NAND3_X2 _10395_ ( .A1(_03074_ ), .A2(fanout_net_13 ), .A3(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ), .ZN(_03230_ ) );
OAI21_X1 _10396_ ( .A(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .B1(_03079_ ), .B2(\u_exu.alu_ctrl[3] ), .ZN(_03231_ ) );
AND3_X4 _10397_ ( .A1(_03229_ ), .A2(_03230_ ), .A3(_03231_ ), .ZN(_03232_ ) );
INV_X1 _10398_ ( .A(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ), .ZN(_03233_ ) );
AND2_X1 _10399_ ( .A1(_03228_ ), .A2(_03233_ ), .ZN(_03234_ ) );
OAI211_X2 _10400_ ( .A(_03222_ ), .B(_03226_ ), .C1(_03232_ ), .C2(_03234_ ), .ZN(_03235_ ) );
AND2_X1 _10401_ ( .A1(_03224_ ), .A2(\u_exu.alu_p1[2] ), .ZN(_03236_ ) );
AND2_X2 _10402_ ( .A1(_03222_ ), .A2(_03236_ ), .ZN(_03237_ ) );
INV_X1 _10403_ ( .A(\u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03238_ ) );
AOI21_X2 _10404_ ( .A(_03237_ ), .B1(_03238_ ), .B2(_03221_ ), .ZN(_03239_ ) );
AOI211_X2 _10405_ ( .A(_03210_ ), .B(_03219_ ), .C1(_03235_ ), .C2(_03239_ ), .ZN(_03240_ ) );
NAND3_X1 _10406_ ( .A1(_03209_ ), .A2(\u_exu.alu_p1[6] ), .A3(_03202_ ), .ZN(_03241_ ) );
INV_X1 _10407_ ( .A(_03208_ ), .ZN(_03242_ ) );
INV_X1 _10408_ ( .A(\u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03243_ ) );
AND2_X1 _10409_ ( .A1(_03216_ ), .A2(_03243_ ), .ZN(_03244_ ) );
AND2_X1 _10410_ ( .A1(_03212_ ), .A2(\u_exu.alu_p1[4] ), .ZN(_03245_ ) );
AOI21_X1 _10411_ ( .A(_03244_ ), .B1(_03217_ ), .B2(_03245_ ), .ZN(_03246_ ) );
OAI221_X4 _10412_ ( .A(_03241_ ), .B1(\u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B2(_03242_ ), .C1(_03246_ ), .C2(_03210_ ), .ZN(_03247_ ) );
NOR2_X2 _10413_ ( .A1(_03240_ ), .A2(_03247_ ), .ZN(_03248_ ) );
INV_X1 _10414_ ( .A(\u_exu.alu_p1[8] ), .ZN(_03249_ ) );
XNOR2_X1 _10415_ ( .A(_03169_ ), .B(_03249_ ), .ZN(_03250_ ) );
NAND3_X1 _10416_ ( .A1(_03177_ ), .A2(_03167_ ), .A3(_03250_ ), .ZN(_03251_ ) );
OR3_X4 _10417_ ( .A1(_03248_ ), .A2(_03189_ ), .A3(_03251_ ), .ZN(_03252_ ) );
AND2_X4 _10418_ ( .A1(_03200_ ), .A2(_03252_ ), .ZN(_03253_ ) );
INV_X4 _10419_ ( .A(_03253_ ), .ZN(_03254_ ) );
NAND2_X2 _10420_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[20] ), .ZN(_03255_ ) );
XNOR2_X1 _10421_ ( .A(_03255_ ), .B(_03141_ ), .ZN(_03256_ ) );
INV_X1 _10422_ ( .A(\u_exu.alu_p1[20] ), .ZN(_03257_ ) );
XNOR2_X1 _10423_ ( .A(_03256_ ), .B(_03257_ ), .ZN(_03258_ ) );
NAND2_X1 _10424_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[21] ), .ZN(_03259_ ) );
XNOR2_X1 _10425_ ( .A(_03259_ ), .B(_03141_ ), .ZN(_03260_ ) );
XNOR2_X1 _10426_ ( .A(_03260_ ), .B(\u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03261_ ) );
AND2_X1 _10427_ ( .A1(_03258_ ), .A2(_03261_ ), .ZN(_03262_ ) );
NAND2_X1 _10428_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[23] ), .ZN(_03263_ ) );
XNOR2_X1 _10429_ ( .A(_03263_ ), .B(_03141_ ), .ZN(_03264_ ) );
INV_X1 _10430_ ( .A(\u_exu.alu_p1[23] ), .ZN(_03265_ ) );
XNOR2_X1 _10431_ ( .A(_03264_ ), .B(_03265_ ), .ZN(_03266_ ) );
NAND2_X2 _10432_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[22] ), .ZN(_03267_ ) );
XNOR2_X2 _10433_ ( .A(_03267_ ), .B(_03142_ ), .ZN(_03268_ ) );
INV_X1 _10434_ ( .A(\u_exu.alu_p1[22] ), .ZN(_03269_ ) );
XNOR2_X1 _10435_ ( .A(_03268_ ), .B(_03269_ ), .ZN(_03270_ ) );
AND3_X1 _10436_ ( .A1(_03262_ ), .A2(_03266_ ), .A3(_03270_ ), .ZN(_03271_ ) );
NAND2_X2 _10437_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[18] ), .ZN(_03272_ ) );
XNOR2_X1 _10438_ ( .A(_03272_ ), .B(_03141_ ), .ZN(_03273_ ) );
INV_X1 _10439_ ( .A(\u_exu.alu_p1[18] ), .ZN(_03274_ ) );
XNOR2_X1 _10440_ ( .A(_03273_ ), .B(_03274_ ), .ZN(_03275_ ) );
NAND2_X4 _10441_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[19] ), .ZN(_03276_ ) );
XNOR2_X2 _10442_ ( .A(_03276_ ), .B(_03141_ ), .ZN(_03277_ ) );
XNOR2_X2 _10443_ ( .A(_03277_ ), .B(\u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03278_ ) );
AND2_X2 _10444_ ( .A1(_03275_ ), .A2(_03278_ ), .ZN(_03279_ ) );
NAND2_X2 _10445_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[16] ), .ZN(_03280_ ) );
XNOR2_X1 _10446_ ( .A(_03280_ ), .B(_03141_ ), .ZN(_03281_ ) );
INV_X1 _10447_ ( .A(\u_exu.alu_p1[16] ), .ZN(_03282_ ) );
XNOR2_X1 _10448_ ( .A(_03281_ ), .B(_03282_ ), .ZN(_03283_ ) );
NAND2_X4 _10449_ ( .A1(_03074_ ), .A2(\u_exu.alu_p2[17] ), .ZN(_03284_ ) );
XNOR2_X2 _10450_ ( .A(_03284_ ), .B(_03141_ ), .ZN(_03285_ ) );
XNOR2_X2 _10451_ ( .A(_03285_ ), .B(\u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03286_ ) );
AND3_X1 _10452_ ( .A1(_03279_ ), .A2(_03283_ ), .A3(_03286_ ), .ZN(_03287_ ) );
NAND3_X4 _10453_ ( .A1(_03254_ ), .A2(_03271_ ), .A3(_03287_ ), .ZN(_03288_ ) );
AND2_X1 _10454_ ( .A1(_03273_ ), .A2(\u_exu.alu_p1[18] ), .ZN(_03289_ ) );
AND2_X1 _10455_ ( .A1(_03278_ ), .A2(_03289_ ), .ZN(_03290_ ) );
INV_X1 _10456_ ( .A(\u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03291_ ) );
AOI21_X1 _10457_ ( .A(_03290_ ), .B1(_03291_ ), .B2(_03277_ ), .ZN(_03292_ ) );
INV_X1 _10458_ ( .A(\u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03293_ ) );
AND2_X1 _10459_ ( .A1(_03285_ ), .A2(_03293_ ), .ZN(_03294_ ) );
AND2_X1 _10460_ ( .A1(_03281_ ), .A2(\u_exu.alu_p1[16] ), .ZN(_03295_ ) );
AOI21_X2 _10461_ ( .A(_03294_ ), .B1(_03286_ ), .B2(_03295_ ), .ZN(_03296_ ) );
INV_X1 _10462_ ( .A(_03296_ ), .ZN(_03297_ ) );
NAND2_X1 _10463_ ( .A1(_03297_ ), .A2(_03279_ ), .ZN(_03298_ ) );
AND2_X2 _10464_ ( .A1(_03292_ ), .A2(_03298_ ), .ZN(_03299_ ) );
AND2_X2 _10465_ ( .A1(_03266_ ), .A2(_03270_ ), .ZN(_03300_ ) );
NAND2_X1 _10466_ ( .A1(_03300_ ), .A2(_03262_ ), .ZN(_03301_ ) );
OR2_X1 _10467_ ( .A1(_03299_ ), .A2(_03301_ ), .ZN(_03302_ ) );
INV_X1 _10468_ ( .A(_03300_ ), .ZN(_03303_ ) );
AND2_X2 _10469_ ( .A1(_03256_ ), .A2(\u_exu.alu_p1[20] ), .ZN(_03304_ ) );
AND2_X1 _10470_ ( .A1(_03261_ ), .A2(_03304_ ), .ZN(_03305_ ) );
INV_X1 _10471_ ( .A(\u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03306_ ) );
AOI21_X1 _10472_ ( .A(_03305_ ), .B1(_03306_ ), .B2(_03260_ ), .ZN(_03307_ ) );
OR2_X1 _10473_ ( .A1(_03303_ ), .A2(_03307_ ), .ZN(_03308_ ) );
AND2_X1 _10474_ ( .A1(_03268_ ), .A2(\u_exu.alu_p1[22] ), .ZN(_03309_ ) );
AND2_X1 _10475_ ( .A1(_03266_ ), .A2(_03309_ ), .ZN(_03310_ ) );
AOI21_X1 _10476_ ( .A(_03310_ ), .B1(\u_exu.alu_p1[23] ), .B2(_03264_ ), .ZN(_03311_ ) );
AND3_X4 _10477_ ( .A1(_03302_ ), .A2(_03308_ ), .A3(_03311_ ), .ZN(_03312_ ) );
AND2_X4 _10478_ ( .A1(_03288_ ), .A2(_03312_ ), .ZN(_03313_ ) );
INV_X4 _10479_ ( .A(_03313_ ), .ZN(_03314_ ) );
NAND2_X1 _10480_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[27] ), .ZN(_03315_ ) );
XNOR2_X1 _10481_ ( .A(_03315_ ), .B(_03142_ ), .ZN(_03316_ ) );
INV_X1 _10482_ ( .A(\u_exu.alu_p1[27] ), .ZN(_03317_ ) );
XNOR2_X1 _10483_ ( .A(_03316_ ), .B(_03317_ ), .ZN(_03318_ ) );
NAND2_X1 _10484_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[26] ), .ZN(_03319_ ) );
XNOR2_X1 _10485_ ( .A(_03319_ ), .B(_03142_ ), .ZN(_03320_ ) );
INV_X1 _10486_ ( .A(\u_exu.alu_p1[26] ), .ZN(_03321_ ) );
XNOR2_X1 _10487_ ( .A(_03320_ ), .B(_03321_ ), .ZN(_03322_ ) );
NAND2_X1 _10488_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[24] ), .ZN(_03323_ ) );
XNOR2_X1 _10489_ ( .A(_03323_ ), .B(_03142_ ), .ZN(_03324_ ) );
INV_X1 _10490_ ( .A(\u_exu.alu_p1[24] ), .ZN(_03325_ ) );
XNOR2_X1 _10491_ ( .A(_03324_ ), .B(_03325_ ), .ZN(_03326_ ) );
NAND2_X1 _10492_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[25] ), .ZN(_03327_ ) );
XNOR2_X1 _10493_ ( .A(_03327_ ), .B(_03142_ ), .ZN(_03328_ ) );
INV_X1 _10494_ ( .A(\u_exu.alu_p1[25] ), .ZN(_03329_ ) );
XNOR2_X1 _10495_ ( .A(_03328_ ), .B(_03329_ ), .ZN(_03330_ ) );
AND2_X1 _10496_ ( .A1(_03326_ ), .A2(_03330_ ), .ZN(_03331_ ) );
NAND4_X4 _10497_ ( .A1(_03314_ ), .A2(_03318_ ), .A3(_03322_ ), .A4(_03331_ ), .ZN(_03332_ ) );
AND2_X1 _10498_ ( .A1(_03324_ ), .A2(\u_exu.alu_p1[24] ), .ZN(_03333_ ) );
AND2_X1 _10499_ ( .A1(_03330_ ), .A2(_03333_ ), .ZN(_03334_ ) );
AOI21_X1 _10500_ ( .A(_03334_ ), .B1(\u_exu.alu_p1[25] ), .B2(_03328_ ), .ZN(_03335_ ) );
INV_X1 _10501_ ( .A(_03318_ ), .ZN(_03336_ ) );
INV_X1 _10502_ ( .A(_03322_ ), .ZN(_03337_ ) );
NOR3_X1 _10503_ ( .A1(_03335_ ), .A2(_03336_ ), .A3(_03337_ ), .ZN(_03338_ ) );
AND2_X1 _10504_ ( .A1(_03316_ ), .A2(\u_exu.alu_p1[27] ), .ZN(_03339_ ) );
AND2_X1 _10505_ ( .A1(_03320_ ), .A2(\u_exu.alu_p1[26] ), .ZN(_03340_ ) );
AND2_X1 _10506_ ( .A1(_03318_ ), .A2(_03340_ ), .ZN(_03341_ ) );
NOR3_X1 _10507_ ( .A1(_03338_ ), .A2(_03339_ ), .A3(_03341_ ), .ZN(_03342_ ) );
AND2_X4 _10508_ ( .A1(_03332_ ), .A2(_03342_ ), .ZN(_03343_ ) );
INV_X4 _10509_ ( .A(_03343_ ), .ZN(_03344_ ) );
NAND2_X1 _10510_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[29] ), .ZN(_03345_ ) );
XNOR2_X1 _10511_ ( .A(_03345_ ), .B(_03142_ ), .ZN(_03346_ ) );
INV_X1 _10512_ ( .A(\u_exu.alu_p1[29] ), .ZN(_03347_ ) );
XNOR2_X1 _10513_ ( .A(_03346_ ), .B(_03347_ ), .ZN(_03348_ ) );
NAND2_X1 _10514_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[28] ), .ZN(_03349_ ) );
XNOR2_X1 _10515_ ( .A(_03349_ ), .B(_03142_ ), .ZN(_03350_ ) );
INV_X1 _10516_ ( .A(\u_exu.alu_p1[28] ), .ZN(_03351_ ) );
XNOR2_X1 _10517_ ( .A(_03350_ ), .B(_03351_ ), .ZN(_03352_ ) );
NAND3_X4 _10518_ ( .A1(_03344_ ), .A2(_03348_ ), .A3(_03352_ ), .ZN(_03353_ ) );
AND2_X1 _10519_ ( .A1(_03350_ ), .A2(\u_exu.alu_p1[28] ), .ZN(_03354_ ) );
AND2_X1 _10520_ ( .A1(_03348_ ), .A2(_03354_ ), .ZN(_03355_ ) );
AOI21_X1 _10521_ ( .A(_03355_ ), .B1(\u_exu.alu_p1[29] ), .B2(_03346_ ), .ZN(_03356_ ) );
AOI21_X4 _10522_ ( .A(_03146_ ), .B1(_03353_ ), .B2(_03356_ ), .ZN(_03357_ ) );
INV_X2 _10523_ ( .A(_03357_ ), .ZN(_03358_ ) );
NAND2_X1 _10524_ ( .A1(_03075_ ), .A2(\u_exu.alu_p2[31] ), .ZN(_03359_ ) );
XNOR2_X1 _10525_ ( .A(_03359_ ), .B(_03142_ ), .ZN(_03360_ ) );
INV_X1 _10526_ ( .A(\u_exu.alu_p1[31] ), .ZN(_03361_ ) );
XNOR2_X1 _10527_ ( .A(_03360_ ), .B(_03361_ ), .ZN(_03362_ ) );
AND2_X1 _10528_ ( .A1(_03143_ ), .A2(\u_exu.alu_p1[30] ), .ZN(_03363_ ) );
INV_X1 _10529_ ( .A(_03363_ ), .ZN(_03364_ ) );
AND3_X4 _10530_ ( .A1(_03358_ ), .A2(_03362_ ), .A3(_03364_ ), .ZN(_03365_ ) );
INV_X1 _10531_ ( .A(\u_exu.alu_ctrl[1] ), .ZN(_03366_ ) );
NOR2_X1 _10532_ ( .A1(_03362_ ), .A2(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ), .ZN(_03367_ ) );
OR3_X4 _10533_ ( .A1(_03365_ ), .A2(_03366_ ), .A3(_03367_ ), .ZN(_03368_ ) );
AND2_X1 _10534_ ( .A1(_03360_ ), .A2(\u_exu.alu_p1[31] ), .ZN(_03369_ ) );
OR2_X1 _10535_ ( .A1(_03369_ ), .A2(_03363_ ), .ZN(_03370_ ) );
OAI221_X1 _10536_ ( .A(_03366_ ), .B1(\u_exu.alu_p1[31] ), .B2(_03360_ ), .C1(_03357_ ), .C2(_03370_ ), .ZN(_03371_ ) );
NAND3_X2 _10537_ ( .A1(_03368_ ), .A2(\u_exu.alu_ctrl[2] ), .A3(_03371_ ), .ZN(_03372_ ) );
INV_X1 _10538_ ( .A(\u_exu.alu_ctrl[5] ), .ZN(_03373_ ) );
NOR2_X1 _10539_ ( .A1(_03373_ ), .A2(\u_exu.alu_ctrl[4] ), .ZN(_03374_ ) );
NAND3_X1 _10540_ ( .A1(_03372_ ), .A2(\u_exu.alu_ctrl[6] ), .A3(_03374_ ), .ZN(_03375_ ) );
AOI21_X1 _10541_ ( .A(\u_exu.alu_ctrl[2] ), .B1(_03368_ ), .B2(_03371_ ), .ZN(_03376_ ) );
OAI21_X1 _10542_ ( .A(_03137_ ), .B1(_03375_ ), .B2(_03376_ ), .ZN(_03377_ ) );
AND2_X2 _10543_ ( .A1(_03069_ ), .A2(\u_exu.alu_ctrl[6] ), .ZN(_03378_ ) );
INV_X2 _10544_ ( .A(fanout_net_20 ), .ZN(_03379_ ) );
AND2_X2 _10545_ ( .A1(_03078_ ), .A2(_03379_ ), .ZN(_03380_ ) );
INV_X1 _10546_ ( .A(_03380_ ), .ZN(_03381_ ) );
NOR2_X1 _10547_ ( .A1(_03274_ ), .A2(fanout_net_13 ), .ZN(_03382_ ) );
AND2_X1 _10548_ ( .A1(\u_exu.alu_p1[19] ), .A2(fanout_net_13 ), .ZN(_03383_ ) );
INV_X1 _10549_ ( .A(fanout_net_15 ), .ZN(_03384_ ) );
OR3_X1 _10550_ ( .A1(_03382_ ), .A2(_03383_ ), .A3(_03384_ ), .ZN(_03385_ ) );
NOR2_X1 _10551_ ( .A1(_03282_ ), .A2(fanout_net_13 ), .ZN(_03386_ ) );
AND2_X1 _10552_ ( .A1(\u_exu.alu_p1[17] ), .A2(fanout_net_13 ), .ZN(_03387_ ) );
OR3_X1 _10553_ ( .A1(_03386_ ), .A2(_03387_ ), .A3(fanout_net_15 ), .ZN(_03388_ ) );
AOI21_X1 _10554_ ( .A(fanout_net_17 ), .B1(_03385_ ), .B2(_03388_ ), .ZN(_03389_ ) );
INV_X1 _10555_ ( .A(fanout_net_17 ), .ZN(_03390_ ) );
NOR2_X1 _10556_ ( .A1(_03257_ ), .A2(fanout_net_13 ), .ZN(_03391_ ) );
AND2_X1 _10557_ ( .A1(\u_exu.alu_p1[21] ), .A2(fanout_net_13 ), .ZN(_03392_ ) );
OR3_X1 _10558_ ( .A1(_03391_ ), .A2(_03392_ ), .A3(fanout_net_15 ), .ZN(_03393_ ) );
AND2_X1 _10559_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1[23] ), .ZN(_03394_ ) );
INV_X1 _10560_ ( .A(_03394_ ), .ZN(_03395_ ) );
OAI211_X1 _10561_ ( .A(_03395_ ), .B(fanout_net_15 ), .C1(fanout_net_13 ), .C2(_03269_ ), .ZN(_03396_ ) );
AOI21_X1 _10562_ ( .A(_03390_ ), .B1(_03393_ ), .B2(_03396_ ), .ZN(_03397_ ) );
NOR2_X1 _10563_ ( .A1(_03389_ ), .A2(_03397_ ), .ZN(_03398_ ) );
NOR2_X1 _10564_ ( .A1(_03321_ ), .A2(fanout_net_13 ), .ZN(_03399_ ) );
AND2_X1 _10565_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1[27] ), .ZN(_03400_ ) );
OR3_X1 _10566_ ( .A1(_03399_ ), .A2(_03400_ ), .A3(_03384_ ), .ZN(_03401_ ) );
NOR2_X1 _10567_ ( .A1(_03325_ ), .A2(fanout_net_13 ), .ZN(_03402_ ) );
INV_X1 _10568_ ( .A(_03402_ ), .ZN(_03403_ ) );
AND2_X1 _10569_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1[25] ), .ZN(_03404_ ) );
INV_X1 _10570_ ( .A(_03404_ ), .ZN(_03405_ ) );
NAND3_X1 _10571_ ( .A1(_03403_ ), .A2(_03384_ ), .A3(_03405_ ), .ZN(_03406_ ) );
AOI21_X1 _10572_ ( .A(fanout_net_17 ), .B1(_03401_ ), .B2(_03406_ ), .ZN(_03407_ ) );
NOR2_X1 _10573_ ( .A1(_03351_ ), .A2(fanout_net_13 ), .ZN(_03408_ ) );
AND2_X1 _10574_ ( .A1(\u_exu.alu_p1[29] ), .A2(fanout_net_13 ), .ZN(_03409_ ) );
OR3_X1 _10575_ ( .A1(_03408_ ), .A2(_03409_ ), .A3(fanout_net_15 ), .ZN(_03410_ ) );
MUX2_X1 _10576_ ( .A(_03144_ ), .B(_03361_ ), .S(fanout_net_13 ), .Z(_03411_ ) );
INV_X1 _10577_ ( .A(_03411_ ), .ZN(_03412_ ) );
BUF_X2 _10578_ ( .A(_03384_ ), .Z(_03413_ ) );
OAI21_X1 _10579_ ( .A(_03410_ ), .B1(_03412_ ), .B2(_03413_ ), .ZN(_03414_ ) );
AOI21_X1 _10580_ ( .A(_03407_ ), .B1(fanout_net_17 ), .B2(_03414_ ), .ZN(_03415_ ) );
MUX2_X1 _10581_ ( .A(_03398_ ), .B(_03415_ ), .S(fanout_net_19 ), .Z(_03416_ ) );
NAND2_X1 _10582_ ( .A1(_03416_ ), .A2(\u_exu.alu_p2[4] ), .ZN(_03417_ ) );
INV_X2 _10583_ ( .A(\u_exu.alu_p2[4] ), .ZN(_03418_ ) );
AND3_X1 _10584_ ( .A1(_03413_ ), .A2(fanout_net_13 ), .A3(\u_exu.alu_p1[1] ), .ZN(_03419_ ) );
AND2_X1 _10585_ ( .A1(_03079_ ), .A2(\u_exu.alu_p1[0] ), .ZN(_03420_ ) );
AND2_X1 _10586_ ( .A1(_03420_ ), .A2(_03384_ ), .ZN(_03421_ ) );
OR2_X1 _10587_ ( .A1(_03421_ ), .A2(fanout_net_17 ), .ZN(_03422_ ) );
MUX2_X1 _10588_ ( .A(\u_exu.alu_p1[2] ), .B(\u_exu.alu_p1[3] ), .S(fanout_net_13 ), .Z(_03423_ ) );
AOI211_X1 _10589_ ( .A(_03419_ ), .B(_03422_ ), .C1(fanout_net_15 ), .C2(_03423_ ), .ZN(_03424_ ) );
NOR2_X1 _10590_ ( .A1(_03203_ ), .A2(fanout_net_13 ), .ZN(_03425_ ) );
AND2_X1 _10591_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1[7] ), .ZN(_03426_ ) );
OR3_X1 _10592_ ( .A1(_03425_ ), .A2(_03426_ ), .A3(_03413_ ), .ZN(_03427_ ) );
NOR2_X1 _10593_ ( .A1(_03213_ ), .A2(fanout_net_13 ), .ZN(_03428_ ) );
AND2_X1 _10594_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1[5] ), .ZN(_03429_ ) );
OR3_X1 _10595_ ( .A1(_03428_ ), .A2(_03429_ ), .A3(fanout_net_15 ), .ZN(_03430_ ) );
NAND2_X1 _10596_ ( .A1(_03427_ ), .A2(_03430_ ), .ZN(_03431_ ) );
AOI211_X1 _10597_ ( .A(fanout_net_19 ), .B(_03424_ ), .C1(fanout_net_17 ), .C2(_03431_ ), .ZN(_03432_ ) );
INV_X1 _10598_ ( .A(fanout_net_19 ), .ZN(_03433_ ) );
NOR2_X1 _10599_ ( .A1(_03184_ ), .A2(fanout_net_13 ), .ZN(_03434_ ) );
AND2_X1 _10600_ ( .A1(\u_exu.alu_p1[13] ), .A2(fanout_net_13 ), .ZN(_03435_ ) );
OAI21_X1 _10601_ ( .A(_03413_ ), .B1(_03434_ ), .B2(_03435_ ), .ZN(_03436_ ) );
NOR2_X1 _10602_ ( .A1(_03179_ ), .A2(fanout_net_13 ), .ZN(_03437_ ) );
AND2_X1 _10603_ ( .A1(\u_exu.alu_p1[15] ), .A2(fanout_net_13 ), .ZN(_03438_ ) );
OAI21_X1 _10604_ ( .A(fanout_net_15 ), .B1(_03437_ ), .B2(_03438_ ), .ZN(_03439_ ) );
NAND2_X1 _10605_ ( .A1(_03436_ ), .A2(_03439_ ), .ZN(_03440_ ) );
NAND2_X1 _10606_ ( .A1(_03440_ ), .A2(fanout_net_17 ), .ZN(_03441_ ) );
NOR2_X1 _10607_ ( .A1(_03175_ ), .A2(fanout_net_13 ), .ZN(_03442_ ) );
AND2_X1 _10608_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[11] ), .ZN(_03443_ ) );
OR3_X1 _10609_ ( .A1(_03442_ ), .A2(_03443_ ), .A3(_03413_ ), .ZN(_03444_ ) );
NOR2_X1 _10610_ ( .A1(_03249_ ), .A2(fanout_net_14 ), .ZN(_03445_ ) );
AND2_X1 _10611_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[9] ), .ZN(_03446_ ) );
OR3_X1 _10612_ ( .A1(_03445_ ), .A2(_03446_ ), .A3(fanout_net_15 ), .ZN(_03447_ ) );
NAND3_X1 _10613_ ( .A1(_03444_ ), .A2(_03447_ ), .A3(_03390_ ), .ZN(_03448_ ) );
AOI21_X1 _10614_ ( .A(_03433_ ), .B1(_03441_ ), .B2(_03448_ ), .ZN(_03449_ ) );
OAI21_X1 _10615_ ( .A(_03418_ ), .B1(_03432_ ), .B2(_03449_ ), .ZN(_03450_ ) );
AOI221_X4 _10616_ ( .A(_03381_ ), .B1(\u_exu.alu_ctrl[1] ), .B2(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_Y_$_MUX__B_A_$_NOR__Y_A_$_ANDNOT__Y_B ), .C1(_03417_ ), .C2(_03450_ ), .ZN(_03451_ ) );
NOR3_X1 _10617_ ( .A1(_03377_ ), .A2(_03378_ ), .A3(_03451_ ), .ZN(_03452_ ) );
BUF_X4 _10618_ ( .A(_03433_ ), .Z(_03453_ ) );
BUF_X4 _10619_ ( .A(_03453_ ), .Z(_03454_ ) );
BUF_X4 _10620_ ( .A(_03390_ ), .Z(_03455_ ) );
BUF_X4 _10621_ ( .A(_03455_ ), .Z(_03456_ ) );
BUF_X4 _10622_ ( .A(_03456_ ), .Z(_03457_ ) );
NAND4_X1 _10623_ ( .A1(_03421_ ), .A2(_03418_ ), .A3(_03454_ ), .A4(_03457_ ), .ZN(_03458_ ) );
AOI211_X1 _10624_ ( .A(_03084_ ), .B(_03452_ ), .C1(_03378_ ), .C2(_03458_ ), .ZN(_03459_ ) );
AND2_X1 _10625_ ( .A1(_03374_ ), .A2(fanout_net_20 ), .ZN(_03460_ ) );
AND2_X1 _10626_ ( .A1(_03110_ ), .A2(_03084_ ), .ZN(_03461_ ) );
NOR3_X2 _10627_ ( .A1(_03459_ ), .A2(_03460_ ), .A3(_03461_ ), .ZN(_03462_ ) );
AND2_X1 _10628_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[0] ), .ZN(_03463_ ) );
INV_X1 _10629_ ( .A(_03463_ ), .ZN(_03464_ ) );
OAI21_X1 _10630_ ( .A(\u_exu.alu_ctrl[0] ), .B1(fanout_net_14 ), .B2(\u_exu.alu_p1[0] ), .ZN(_03465_ ) );
AND3_X1 _10631_ ( .A1(_03460_ ), .A2(_03464_ ), .A3(_03465_ ), .ZN(_03466_ ) );
OAI221_X2 _10632_ ( .A(_03071_ ), .B1(_03076_ ), .B2(_03082_ ), .C1(_03462_ ), .C2(_03466_ ), .ZN(_03467_ ) );
NAND4_X1 _10633_ ( .A1(_03373_ ), .A2(_03077_ ), .A3(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ), .A4(fanout_net_20 ), .ZN(_03468_ ) );
AND3_X4 _10634_ ( .A1(_03467_ ), .A2(_01450_ ), .A3(_03468_ ), .ZN(_03469_ ) );
BUF_X4 _10635_ ( .A(_00747_ ), .Z(_03470_ ) );
INV_X2 _10636_ ( .A(_03470_ ), .ZN(_03471_ ) );
NOR2_X4 _10637_ ( .A1(_03469_ ), .A2(_03471_ ), .ZN(_03472_ ) );
BUF_X8 _10638_ ( .A(_03472_ ), .Z(_03473_ ) );
NAND3_X1 _10639_ ( .A1(_01053_ ), .A2(_00895_ ), .A3(_01480_ ), .ZN(_03474_ ) );
BUF_X4 _10640_ ( .A(_03474_ ), .Z(_03475_ ) );
NOR2_X1 _10641_ ( .A1(_01459_ ), .A2(_01565_ ), .ZN(_03476_ ) );
INV_X1 _10642_ ( .A(_03476_ ), .ZN(_03477_ ) );
BUF_X4 _10643_ ( .A(_03477_ ), .Z(_03478_ ) );
AND3_X1 _10644_ ( .A1(_01422_ ), .A2(_01418_ ), .A3(_01445_ ), .ZN(_03479_ ) );
NOR2_X1 _10645_ ( .A1(_00694_ ), .A2(_00741_ ), .ZN(_03480_ ) );
AND2_X2 _10646_ ( .A1(_00669_ ), .A2(_03480_ ), .ZN(_03481_ ) );
BUF_X4 _10647_ ( .A(_03481_ ), .Z(_03482_ ) );
BUF_X2 _10648_ ( .A(_00919_ ), .Z(_03483_ ) );
XNOR2_X1 _10649_ ( .A(_03483_ ), .B(_01235_ ), .ZN(_03484_ ) );
XNOR2_X1 _10650_ ( .A(_00955_ ), .B(_01226_ ), .ZN(_03485_ ) );
XNOR2_X1 _10651_ ( .A(_01044_ ), .B(_01230_ ), .ZN(_03486_ ) );
BUF_X4 _10652_ ( .A(_00921_ ), .Z(_03487_ ) );
XNOR2_X1 _10653_ ( .A(_03487_ ), .B(_01239_ ), .ZN(_03488_ ) );
AND4_X1 _10654_ ( .A1(_03484_ ), .A2(_03485_ ), .A3(_03486_ ), .A4(_03488_ ), .ZN(_03489_ ) );
AND2_X1 _10655_ ( .A1(_01223_ ), .A2(_03489_ ), .ZN(_03490_ ) );
INV_X1 _10656_ ( .A(_03490_ ), .ZN(_03491_ ) );
BUF_X2 _10657_ ( .A(_03491_ ), .Z(_03492_ ) );
BUF_X2 _10658_ ( .A(_00971_ ), .Z(_03493_ ) );
BUF_X4 _10659_ ( .A(_00955_ ), .Z(_03494_ ) );
NAND3_X1 _10660_ ( .A1(_03494_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03495_ ) );
NAND2_X1 _10661_ ( .A1(_03495_ ), .A2(_03487_ ), .ZN(_03496_ ) );
BUF_X2 _10662_ ( .A(_03483_ ), .Z(_03497_ ) );
BUF_X2 _10663_ ( .A(_00875_ ), .Z(_03498_ ) );
NAND3_X1 _10664_ ( .A1(_03497_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03499_ ) );
NAND3_X1 _10665_ ( .A1(_03497_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03500_ ) );
NAND2_X1 _10666_ ( .A1(_03499_ ), .A2(_03500_ ), .ZN(_03501_ ) );
BUF_X4 _10667_ ( .A(_00988_ ), .Z(_03502_ ) );
BUF_X4 _10668_ ( .A(_03502_ ), .Z(_03503_ ) );
AOI211_X1 _10669_ ( .A(_03496_ ), .B(_03501_ ), .C1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03503_ ), .ZN(_03504_ ) );
BUF_X4 _10670_ ( .A(_03487_ ), .Z(_03505_ ) );
BUF_X4 _10671_ ( .A(_00996_ ), .Z(_03506_ ) );
BUF_X4 _10672_ ( .A(_03506_ ), .Z(_03507_ ) );
AOI21_X1 _10673_ ( .A(_03505_ ), .B1(_03507_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03508_ ) );
BUF_X4 _10674_ ( .A(_03483_ ), .Z(_03509_ ) );
AND3_X1 _10675_ ( .A1(_03509_ ), .A2(_00875_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03510_ ) );
AND2_X1 _10676_ ( .A1(_03483_ ), .A2(fanout_net_22 ), .ZN(_03511_ ) );
BUF_X4 _10677_ ( .A(_03511_ ), .Z(_03512_ ) );
AOI221_X4 _10678_ ( .A(_03510_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03502_ ), .ZN(_03513_ ) );
AOI211_X1 _10679_ ( .A(_03493_ ), .B(_03504_ ), .C1(_03508_ ), .C2(_03513_ ), .ZN(_03514_ ) );
BUF_X4 _10680_ ( .A(_03494_ ), .Z(_03515_ ) );
AND3_X1 _10681_ ( .A1(_03515_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03516_ ) );
BUF_X4 _10682_ ( .A(_00972_ ), .Z(_03517_ ) );
AND2_X1 _10683_ ( .A1(_03494_ ), .A2(\u_reg.rf[1][31] ), .ZN(_03518_ ) );
BUF_X2 _10684_ ( .A(_03509_ ), .Z(_03519_ ) );
OAI21_X1 _10685_ ( .A(_03517_ ), .B1(_03518_ ), .B2(_03519_ ), .ZN(_03520_ ) );
BUF_X4 _10686_ ( .A(_00920_ ), .Z(_03521_ ) );
BUF_X4 _10687_ ( .A(_03521_ ), .Z(_03522_ ) );
AOI211_X1 _10688_ ( .A(_03516_ ), .B(_03520_ ), .C1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03522_ ), .ZN(_03523_ ) );
BUF_X4 _10689_ ( .A(_03517_ ), .Z(_03524_ ) );
BUF_X4 _10690_ ( .A(_03509_ ), .Z(_03525_ ) );
NAND3_X1 _10691_ ( .A1(_03525_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03526_ ) );
NAND3_X1 _10692_ ( .A1(_03515_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03527_ ) );
NAND3_X1 _10693_ ( .A1(_03494_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03528_ ) );
NAND3_X1 _10694_ ( .A1(_03526_ ), .A2(_03527_ ), .A3(_03528_ ), .ZN(_03529_ ) );
BUF_X4 _10695_ ( .A(_03502_ ), .Z(_03530_ ) );
BUF_X4 _10696_ ( .A(_03530_ ), .Z(_03531_ ) );
AOI211_X1 _10697_ ( .A(_03524_ ), .B(_03529_ ), .C1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03531_ ), .ZN(_03532_ ) );
NOR3_X1 _10698_ ( .A1(_03523_ ), .A2(_03532_ ), .A3(_01044_ ), .ZN(_03533_ ) );
OR2_X1 _10699_ ( .A1(_03514_ ), .A2(_03533_ ), .ZN(_03534_ ) );
AOI21_X1 _10700_ ( .A(_03482_ ), .B1(_03492_ ), .B2(_03534_ ), .ZN(_03535_ ) );
AND2_X1 _10701_ ( .A1(_01297_ ), .A2(_01301_ ), .ZN(\ar_data[31] ) );
BUF_X4 _10702_ ( .A(_03491_ ), .Z(_03536_ ) );
BUF_X4 _10703_ ( .A(_03536_ ), .Z(_03537_ ) );
OAI21_X1 _10704_ ( .A(_03535_ ), .B1(\ar_data[31] ), .B2(_03537_ ), .ZN(_03538_ ) );
INV_X1 _10705_ ( .A(_01418_ ), .ZN(_03539_ ) );
BUF_X4 _10706_ ( .A(_03539_ ), .Z(_03540_ ) );
BUF_X4 _10707_ ( .A(_03540_ ), .Z(_03541_ ) );
AOI211_X1 _10708_ ( .A(_03478_ ), .B(_03479_ ), .C1(_03538_ ), .C2(_03541_ ), .ZN(_03542_ ) );
AOI21_X1 _10709_ ( .A(_03542_ ), .B1(_01861_ ), .B2(_01480_ ), .ZN(_03543_ ) );
OAI22_X1 _10710_ ( .A1(_03473_ ), .A2(_03475_ ), .B1(_01805_ ), .B2(_03543_ ), .ZN(_00161_ ) );
NOR2_X1 _10711_ ( .A1(_01564_ ), .A2(_02407_ ), .ZN(_03544_ ) );
BUF_X4 _10712_ ( .A(_03477_ ), .Z(_03545_ ) );
BUF_X4 _10713_ ( .A(_03490_ ), .Z(_03546_ ) );
AOI21_X1 _10714_ ( .A(_03482_ ), .B1(_01530_ ), .B2(_03546_ ), .ZN(_03547_ ) );
BUF_X4 _10715_ ( .A(_03546_ ), .Z(_03548_ ) );
BUF_X4 _10716_ ( .A(_03512_ ), .Z(_03549_ ) );
AOI22_X1 _10717_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03550_ ) );
BUF_X4 _10718_ ( .A(_03530_ ), .Z(_03551_ ) );
AOI22_X1 _10719_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03507_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03552_ ) );
BUF_X2 _10720_ ( .A(_03524_ ), .Z(_03553_ ) );
NAND3_X1 _10721_ ( .A1(_03550_ ), .A2(_03552_ ), .A3(_03553_ ), .ZN(_03554_ ) );
AOI22_X1 _10722_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03555_ ) );
AOI22_X1 _10723_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03507_ ), .B1(_03531_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03556_ ) );
BUF_X4 _10724_ ( .A(_03505_ ), .Z(_03557_ ) );
NAND3_X1 _10725_ ( .A1(_03555_ ), .A2(_03556_ ), .A3(_03557_ ), .ZN(_03558_ ) );
BUF_X2 _10726_ ( .A(_01044_ ), .Z(_03559_ ) );
AND3_X1 _10727_ ( .A1(_03554_ ), .A2(_03558_ ), .A3(_03559_ ), .ZN(_03560_ ) );
BUF_X2 _10728_ ( .A(_03493_ ), .Z(_03561_ ) );
BUF_X4 _10729_ ( .A(_00996_ ), .Z(_03562_ ) );
BUF_X4 _10730_ ( .A(_03562_ ), .Z(_03563_ ) );
AND2_X1 _10731_ ( .A1(_00955_ ), .A2(fanout_net_23 ), .ZN(_03564_ ) );
BUF_X4 _10732_ ( .A(_03564_ ), .Z(_03565_ ) );
BUF_X4 _10733_ ( .A(_03565_ ), .Z(_03566_ ) );
AOI22_X1 _10734_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03567_ ) );
BUF_X4 _10735_ ( .A(_03521_ ), .Z(_03568_ ) );
AOI22_X1 _10736_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03569_ ) );
BUF_X4 _10737_ ( .A(_03487_ ), .Z(_03570_ ) );
BUF_X2 _10738_ ( .A(_03570_ ), .Z(_03571_ ) );
NAND3_X1 _10739_ ( .A1(_03567_ ), .A2(_03569_ ), .A3(_03571_ ), .ZN(_03572_ ) );
BUF_X4 _10740_ ( .A(_00980_ ), .Z(_03573_ ) );
BUF_X4 _10741_ ( .A(_00981_ ), .Z(_03574_ ) );
OAI21_X1 _10742_ ( .A(_03573_ ), .B1(_03574_ ), .B2(_01507_ ), .ZN(_03575_ ) );
BUF_X4 _10743_ ( .A(_03525_ ), .Z(_03576_ ) );
BUF_X4 _10744_ ( .A(_03576_ ), .Z(_03577_ ) );
BUF_X2 _10745_ ( .A(_00875_ ), .Z(_03578_ ) );
BUF_X2 _10746_ ( .A(_03578_ ), .Z(_03579_ ) );
NAND3_X1 _10747_ ( .A1(_03577_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03580_ ) );
BUF_X4 _10748_ ( .A(_03525_ ), .Z(_03581_ ) );
BUF_X4 _10749_ ( .A(_03581_ ), .Z(_03582_ ) );
NAND3_X1 _10750_ ( .A1(_03582_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03583_ ) );
NAND4_X1 _10751_ ( .A1(_03575_ ), .A2(_03553_ ), .A3(_03580_ ), .A4(_03583_ ), .ZN(_03584_ ) );
AND2_X1 _10752_ ( .A1(_03572_ ), .A2(_03584_ ), .ZN(_03585_ ) );
AOI21_X1 _10753_ ( .A(_03560_ ), .B1(_03561_ ), .B2(_03585_ ), .ZN(_03586_ ) );
OAI21_X1 _10754_ ( .A(_03547_ ), .B1(_03548_ ), .B2(_03586_ ), .ZN(_03587_ ) );
AOI21_X1 _10755_ ( .A(_03545_ ), .B1(_03587_ ), .B2(_03541_ ), .ZN(_03588_ ) );
BUF_X4 _10756_ ( .A(_01418_ ), .Z(_03589_ ) );
NAND3_X1 _10757_ ( .A1(_01536_ ), .A2(_03589_ ), .A3(_01552_ ), .ZN(_03590_ ) );
AOI21_X1 _10758_ ( .A(_03544_ ), .B1(_03588_ ), .B2(_03590_ ), .ZN(_03591_ ) );
OAI22_X1 _10759_ ( .A1(_03473_ ), .A2(_03475_ ), .B1(_01805_ ), .B2(_03591_ ), .ZN(_00162_ ) );
BUF_X4 _10760_ ( .A(_01804_ ), .Z(_03592_ ) );
NOR3_X1 _10761_ ( .A1(_01633_ ), .A2(_03540_ ), .A3(_01634_ ), .ZN(_03593_ ) );
BUF_X4 _10762_ ( .A(_03481_ ), .Z(_03594_ ) );
AOI21_X1 _10763_ ( .A(_03594_ ), .B1(_01614_ ), .B2(_03548_ ), .ZN(_03595_ ) );
BUF_X2 _10764_ ( .A(_03524_ ), .Z(_03596_ ) );
AOI22_X1 _10765_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03507_ ), .B1(_03531_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03597_ ) );
NAND3_X1 _10766_ ( .A1(_03582_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03598_ ) );
BUF_X4 _10767_ ( .A(_03494_ ), .Z(_03599_ ) );
BUF_X2 _10768_ ( .A(_03599_ ), .Z(_03600_ ) );
NAND3_X1 _10769_ ( .A1(_03600_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03601_ ) );
AND4_X1 _10770_ ( .A1(_03596_ ), .A2(_03597_ ), .A3(_03598_ ), .A4(_03601_ ), .ZN(_03602_ ) );
BUF_X4 _10771_ ( .A(_03515_ ), .Z(_03603_ ) );
NAND3_X1 _10772_ ( .A1(_03603_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03604_ ) );
NAND2_X1 _10773_ ( .A1(_03604_ ), .A2(_03570_ ), .ZN(_03605_ ) );
BUF_X4 _10774_ ( .A(_03509_ ), .Z(_03606_ ) );
BUF_X4 _10775_ ( .A(_03606_ ), .Z(_03607_ ) );
NAND3_X1 _10776_ ( .A1(_03607_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03608_ ) );
BUF_X4 _10777_ ( .A(_03606_ ), .Z(_03609_ ) );
NAND3_X1 _10778_ ( .A1(_03609_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03610_ ) );
NAND2_X1 _10779_ ( .A1(_03608_ ), .A2(_03610_ ), .ZN(_03611_ ) );
BUF_X4 _10780_ ( .A(_03551_ ), .Z(_03612_ ) );
AOI211_X1 _10781_ ( .A(_03605_ ), .B(_03611_ ), .C1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03612_ ), .ZN(_03613_ ) );
BUF_X2 _10782_ ( .A(_03493_ ), .Z(_03614_ ) );
NOR3_X1 _10783_ ( .A1(_03602_ ), .A2(_03613_ ), .A3(_03614_ ), .ZN(_03615_ ) );
BUF_X4 _10784_ ( .A(_00996_ ), .Z(_03616_ ) );
BUF_X4 _10785_ ( .A(_03616_ ), .Z(_03617_ ) );
BUF_X4 _10786_ ( .A(_03565_ ), .Z(_03618_ ) );
BUF_X4 _10787_ ( .A(_03618_ ), .Z(_03619_ ) );
AOI22_X1 _10788_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03620_ ) );
BUF_X4 _10789_ ( .A(_03517_ ), .Z(_03621_ ) );
BUF_X4 _10790_ ( .A(_03621_ ), .Z(_03622_ ) );
AOI21_X1 _10791_ ( .A(_03622_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03623_ ) );
BUF_X4 _10792_ ( .A(_03582_ ), .Z(_03624_ ) );
NAND3_X1 _10793_ ( .A1(_03624_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03625_ ) );
NAND3_X1 _10794_ ( .A1(_03620_ ), .A2(_03623_ ), .A3(_03625_ ), .ZN(_03626_ ) );
BUF_X4 _10795_ ( .A(_03599_ ), .Z(_03627_ ) );
NAND3_X1 _10796_ ( .A1(_03627_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03628_ ) );
BUF_X4 _10797_ ( .A(_00876_ ), .Z(_03629_ ) );
NAND3_X1 _10798_ ( .A1(_03576_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03630_ ) );
NAND2_X1 _10799_ ( .A1(_03628_ ), .A2(_03630_ ), .ZN(_03631_ ) );
BUF_X2 _10800_ ( .A(_03505_ ), .Z(_03632_ ) );
AOI21_X1 _10801_ ( .A(_03576_ ), .B1(\u_reg.rf[1][21] ), .B2(_03627_ ), .ZN(_03633_ ) );
OR3_X1 _10802_ ( .A1(_03631_ ), .A2(_03632_ ), .A3(_03633_ ), .ZN(_03634_ ) );
AND2_X1 _10803_ ( .A1(_03634_ ), .A2(_03561_ ), .ZN(_03635_ ) );
AOI21_X1 _10804_ ( .A(_03615_ ), .B1(_03626_ ), .B2(_03635_ ), .ZN(_03636_ ) );
OAI21_X1 _10805_ ( .A(_03595_ ), .B1(_03548_ ), .B2(_03636_ ), .ZN(_03637_ ) );
BUF_X4 _10806_ ( .A(_03540_ ), .Z(_03638_ ) );
BUF_X4 _10807_ ( .A(_03638_ ), .Z(_03639_ ) );
AOI211_X1 _10808_ ( .A(_03478_ ), .B(_03593_ ), .C1(_03637_ ), .C2(_03639_ ), .ZN(_03640_ ) );
AND2_X1 _10809_ ( .A1(_01642_ ), .A2(_01861_ ), .ZN(_03641_ ) );
OAI21_X1 _10810_ ( .A(_03592_ ), .B1(_03640_ ), .B2(_03641_ ), .ZN(_03642_ ) );
OAI21_X1 _10811_ ( .A(_03642_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00163_ ) );
CLKBUF_X2 _10812_ ( .A(_01418_ ), .Z(_03643_ ) );
AND3_X1 _10813_ ( .A1(_01696_ ), .A2(_03643_ ), .A3(_01714_ ), .ZN(_03644_ ) );
AOI21_X1 _10814_ ( .A(_03594_ ), .B1(_01688_ ), .B2(_03548_ ), .ZN(_03645_ ) );
BUF_X2 _10815_ ( .A(_03487_ ), .Z(_03646_ ) );
BUF_X4 _10816_ ( .A(_03502_ ), .Z(_03647_ ) );
BUF_X4 _10817_ ( .A(_03647_ ), .Z(_03648_ ) );
AOI21_X1 _10818_ ( .A(_03646_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03649_ ) );
BUF_X4 _10819_ ( .A(_03494_ ), .Z(_03650_ ) );
BUF_X2 _10820_ ( .A(_03650_ ), .Z(_03651_ ) );
BUF_X4 _10821_ ( .A(_01639_ ), .Z(_03652_ ) );
NAND3_X1 _10822_ ( .A1(_03651_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03653_ ) );
NAND3_X1 _10823_ ( .A1(_03582_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03654_ ) );
NAND3_X1 _10824_ ( .A1(_03651_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03655_ ) );
NAND4_X1 _10825_ ( .A1(_03649_ ), .A2(_03653_ ), .A3(_03654_ ), .A4(_03655_ ), .ZN(_03656_ ) );
AOI21_X1 _10826_ ( .A(_03621_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03657_ ) );
NAND3_X1 _10827_ ( .A1(_03651_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03658_ ) );
NAND3_X1 _10828_ ( .A1(_03582_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03659_ ) );
NAND3_X1 _10829_ ( .A1(_03600_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03660_ ) );
NAND4_X1 _10830_ ( .A1(_03657_ ), .A2(_03658_ ), .A3(_03659_ ), .A4(_03660_ ), .ZN(_03661_ ) );
BUF_X2 _10831_ ( .A(_01044_ ), .Z(_03662_ ) );
AND3_X1 _10832_ ( .A1(_03656_ ), .A2(_03661_ ), .A3(_03662_ ), .ZN(_03663_ ) );
OAI21_X1 _10833_ ( .A(_03573_ ), .B1(_03574_ ), .B2(_01653_ ), .ZN(_03664_ ) );
NAND3_X1 _10834_ ( .A1(_03624_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03665_ ) );
NAND3_X1 _10835_ ( .A1(_03624_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03666_ ) );
NAND4_X1 _10836_ ( .A1(_03664_ ), .A2(_03622_ ), .A3(_03665_ ), .A4(_03666_ ), .ZN(_03667_ ) );
AOI22_X1 _10837_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03668_ ) );
AOI22_X1 _10838_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03669_ ) );
NAND3_X1 _10839_ ( .A1(_03668_ ), .A2(_03669_ ), .A3(_03571_ ), .ZN(_03670_ ) );
AND2_X1 _10840_ ( .A1(_03670_ ), .A2(_03561_ ), .ZN(_03671_ ) );
AOI21_X1 _10841_ ( .A(_03663_ ), .B1(_03667_ ), .B2(_03671_ ), .ZN(_03672_ ) );
OAI21_X1 _10842_ ( .A(_03645_ ), .B1(_03548_ ), .B2(_03672_ ), .ZN(_03673_ ) );
AOI211_X1 _10843_ ( .A(_03478_ ), .B(_03644_ ), .C1(_03673_ ), .C2(_03639_ ), .ZN(_03674_ ) );
AND2_X1 _10844_ ( .A1(_01718_ ), .A2(_01861_ ), .ZN(_03675_ ) );
OAI21_X1 _10845_ ( .A(_03592_ ), .B1(_03674_ ), .B2(_03675_ ), .ZN(_03676_ ) );
OAI21_X1 _10846_ ( .A(_03676_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00164_ ) );
AND2_X4 _10847_ ( .A1(_03469_ ), .A2(_01480_ ), .ZN(_03677_ ) );
NOR2_X1 _10848_ ( .A1(_01801_ ), .A2(_03470_ ), .ZN(_03678_ ) );
OAI21_X2 _10849_ ( .A(_01054_ ), .B1(_03677_ ), .B2(_03678_ ), .ZN(_03679_ ) );
NOR2_X1 _10850_ ( .A1(\ar_data[19] ), .A2(_03492_ ), .ZN(_03680_ ) );
INV_X1 _10851_ ( .A(_03481_ ), .ZN(_03681_ ) );
AND3_X1 _10852_ ( .A1(_03483_ ), .A2(_00751_ ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03682_ ) );
AOI221_X4 _10853_ ( .A(_03682_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03502_ ), .ZN(_03683_ ) );
BUF_X4 _10854_ ( .A(_03515_ ), .Z(_03684_ ) );
NAND3_X1 _10855_ ( .A1(_03684_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03685_ ) );
NAND3_X1 _10856_ ( .A1(_03683_ ), .A2(_03570_ ), .A3(_03685_ ), .ZN(_03686_ ) );
AOI22_X1 _10857_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03506_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03687_ ) );
BUF_X2 _10858_ ( .A(_03497_ ), .Z(_03688_ ) );
BUF_X2 _10859_ ( .A(_03498_ ), .Z(_03689_ ) );
NAND3_X1 _10860_ ( .A1(_03688_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03690_ ) );
NAND3_X1 _10861_ ( .A1(_03688_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03691_ ) );
NAND4_X1 _10862_ ( .A1(_03687_ ), .A2(_03621_ ), .A3(_03690_ ), .A4(_03691_ ), .ZN(_03692_ ) );
AND3_X1 _10863_ ( .A1(_03686_ ), .A2(_01044_ ), .A3(_03692_ ), .ZN(_03693_ ) );
AOI22_X1 _10864_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03694_ ) );
BUF_X4 _10865_ ( .A(_03531_ ), .Z(_03695_ ) );
AOI21_X1 _10866_ ( .A(_03596_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03696_ ) );
BUF_X4 _10867_ ( .A(_03609_ ), .Z(_03697_ ) );
BUF_X4 _10868_ ( .A(_03629_ ), .Z(_03698_ ) );
NAND3_X1 _10869_ ( .A1(_03697_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03699_ ) );
NAND3_X1 _10870_ ( .A1(_03694_ ), .A2(_03696_ ), .A3(_03699_ ), .ZN(_03700_ ) );
AOI22_X1 _10871_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03701_ ) );
BUF_X4 _10872_ ( .A(_03524_ ), .Z(_03702_ ) );
OAI21_X1 _10873_ ( .A(_00980_ ), .B1(_03574_ ), .B2(_01751_ ), .ZN(_03703_ ) );
NAND3_X1 _10874_ ( .A1(_03701_ ), .A2(_03702_ ), .A3(_03703_ ), .ZN(_03704_ ) );
BUF_X2 _10875_ ( .A(_03493_ ), .Z(_03705_ ) );
AND2_X1 _10876_ ( .A1(_03704_ ), .A2(_03705_ ), .ZN(_03706_ ) );
AOI21_X1 _10877_ ( .A(_03693_ ), .B1(_03700_ ), .B2(_03706_ ), .ZN(_03707_ ) );
OAI21_X1 _10878_ ( .A(_03681_ ), .B1(_03546_ ), .B2(_03707_ ), .ZN(_03708_ ) );
OAI21_X1 _10879_ ( .A(_03638_ ), .B1(_03680_ ), .B2(_03708_ ), .ZN(_03709_ ) );
NAND3_X1 _10880_ ( .A1(_01774_ ), .A2(_01789_ ), .A3(_03643_ ), .ZN(_03710_ ) );
AND3_X1 _10881_ ( .A1(_03709_ ), .A2(_03476_ ), .A3(_03710_ ), .ZN(_03711_ ) );
BUF_X4 _10882_ ( .A(_01465_ ), .Z(_03712_ ) );
BUF_X4 _10883_ ( .A(_01081_ ), .Z(_03713_ ) );
AOI21_X1 _10884_ ( .A(_01801_ ), .B1(_03712_ ), .B2(_03713_ ), .ZN(_03714_ ) );
OAI21_X1 _10885_ ( .A(_01078_ ), .B1(_03711_ ), .B2(_03714_ ), .ZN(_03715_ ) );
AOI21_X1 _10886_ ( .A(_01076_ ), .B1(_03679_ ), .B2(_03715_ ), .ZN(_00165_ ) );
NOR2_X1 _10887_ ( .A1(_01866_ ), .A2(_03470_ ), .ZN(_03716_ ) );
OAI21_X2 _10888_ ( .A(_01054_ ), .B1(_03677_ ), .B2(_03716_ ), .ZN(_03717_ ) );
NOR2_X1 _10889_ ( .A1(\ar_data[18] ), .A2(_03492_ ), .ZN(_03718_ ) );
AOI21_X1 _10890_ ( .A(_03487_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03719_ ) );
NAND3_X1 _10891_ ( .A1(_03684_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03720_ ) );
BUF_X2 _10892_ ( .A(_03497_ ), .Z(_03721_ ) );
BUF_X2 _10893_ ( .A(_03498_ ), .Z(_03722_ ) );
NAND3_X1 _10894_ ( .A1(_03721_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03723_ ) );
NAND3_X1 _10895_ ( .A1(_03684_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03724_ ) );
NAND4_X1 _10896_ ( .A1(_03719_ ), .A2(_03720_ ), .A3(_03723_ ), .A4(_03724_ ), .ZN(_03725_ ) );
AOI21_X1 _10897_ ( .A(_03517_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03726_ ) );
NAND3_X1 _10898_ ( .A1(_03581_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03727_ ) );
NAND3_X1 _10899_ ( .A1(_03684_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03728_ ) );
NAND3_X1 _10900_ ( .A1(_03684_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03729_ ) );
NAND4_X1 _10901_ ( .A1(_03726_ ), .A2(_03727_ ), .A3(_03728_ ), .A4(_03729_ ), .ZN(_03730_ ) );
AND3_X1 _10902_ ( .A1(_03725_ ), .A2(_03730_ ), .A3(_01044_ ), .ZN(_03731_ ) );
AND3_X1 _10903_ ( .A1(_03519_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03732_ ) );
AND3_X1 _10904_ ( .A1(_03606_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03733_ ) );
BUF_X2 _10905_ ( .A(_03497_ ), .Z(_03734_ ) );
AOI21_X1 _10906_ ( .A(_03734_ ), .B1(\u_reg.rf[1][18] ), .B2(_03650_ ), .ZN(_03735_ ) );
OR4_X1 _10907_ ( .A1(_03646_ ), .A2(_03732_ ), .A3(_03733_ ), .A4(_03735_ ), .ZN(_03736_ ) );
AOI22_X1 _10908_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03565_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03737_ ) );
AOI22_X1 _10909_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03738_ ) );
NAND3_X1 _10910_ ( .A1(_03737_ ), .A2(_03738_ ), .A3(_03646_ ), .ZN(_03739_ ) );
AND2_X1 _10911_ ( .A1(_03739_ ), .A2(_03705_ ), .ZN(_03740_ ) );
AOI21_X1 _10912_ ( .A(_03731_ ), .B1(_03736_ ), .B2(_03740_ ), .ZN(_03741_ ) );
OAI21_X1 _10913_ ( .A(_03681_ ), .B1(_03546_ ), .B2(_03741_ ), .ZN(_03742_ ) );
OAI21_X1 _10914_ ( .A(_03638_ ), .B1(_03718_ ), .B2(_03742_ ), .ZN(_03743_ ) );
NAND3_X1 _10915_ ( .A1(_01871_ ), .A2(_03643_ ), .A3(_01878_ ), .ZN(_03744_ ) );
AND3_X1 _10916_ ( .A1(_03743_ ), .A2(_03476_ ), .A3(_03744_ ), .ZN(_03745_ ) );
BUF_X4 _10917_ ( .A(_02407_ ), .Z(_03746_ ) );
NOR2_X1 _10918_ ( .A1(_01866_ ), .A2(_03746_ ), .ZN(_03747_ ) );
OAI21_X1 _10919_ ( .A(_01078_ ), .B1(_03745_ ), .B2(_03747_ ), .ZN(_03748_ ) );
AOI21_X1 _10920_ ( .A(_01076_ ), .B1(_03717_ ), .B2(_03748_ ), .ZN(_00166_ ) );
NOR2_X1 _10921_ ( .A1(_01940_ ), .A2(_03470_ ), .ZN(_03749_ ) );
OAI21_X2 _10922_ ( .A(_01054_ ), .B1(_03677_ ), .B2(_03749_ ), .ZN(_03750_ ) );
AOI22_X1 _10923_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03751_ ) );
BUF_X2 _10924_ ( .A(_03525_ ), .Z(_03752_ ) );
NAND3_X1 _10925_ ( .A1(_03752_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03753_ ) );
NAND3_X1 _10926_ ( .A1(_03607_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03754_ ) );
NAND4_X1 _10927_ ( .A1(_03751_ ), .A2(_03702_ ), .A3(_03753_ ), .A4(_03754_ ), .ZN(_03755_ ) );
AOI21_X1 _10928_ ( .A(_03524_ ), .B1(_03531_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03756_ ) );
NAND3_X1 _10929_ ( .A1(_03607_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03757_ ) );
NAND3_X1 _10930_ ( .A1(_03627_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03758_ ) );
NAND3_X1 _10931_ ( .A1(_03603_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03759_ ) );
NAND4_X1 _10932_ ( .A1(_03756_ ), .A2(_03757_ ), .A3(_03758_ ), .A4(_03759_ ), .ZN(_03760_ ) );
NAND3_X1 _10933_ ( .A1(_03755_ ), .A2(_03559_ ), .A3(_03760_ ), .ZN(_03761_ ) );
AOI22_X1 _10934_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03507_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03762_ ) );
AOI22_X1 _10935_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03763_ ) );
NAND3_X1 _10936_ ( .A1(_03762_ ), .A2(_03763_ ), .A3(_03557_ ), .ZN(_03764_ ) );
NAND2_X1 _10937_ ( .A1(_03764_ ), .A2(_03614_ ), .ZN(_03765_ ) );
AND3_X1 _10938_ ( .A1(_03609_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03766_ ) );
AND3_X1 _10939_ ( .A1(_03721_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03767_ ) );
AOI21_X1 _10940_ ( .A(_03576_ ), .B1(\u_reg.rf[1][17] ), .B2(_03603_ ), .ZN(_03768_ ) );
NOR4_X1 _10941_ ( .A1(_03766_ ), .A2(_03767_ ), .A3(_03768_ ), .A4(_03646_ ), .ZN(_03769_ ) );
OAI21_X1 _10942_ ( .A(_03761_ ), .B1(_03765_ ), .B2(_03769_ ), .ZN(_03770_ ) );
AOI21_X1 _10943_ ( .A(_03482_ ), .B1(_03536_ ), .B2(_03770_ ), .ZN(_03771_ ) );
OAI21_X1 _10944_ ( .A(_03771_ ), .B1(\ar_data[17] ), .B2(_03492_ ), .ZN(_03772_ ) );
AOI21_X1 _10945_ ( .A(_03477_ ), .B1(_03772_ ), .B2(_03638_ ), .ZN(_03773_ ) );
NAND3_X1 _10946_ ( .A1(_01932_ ), .A2(_03589_ ), .A3(_01933_ ), .ZN(_03774_ ) );
AND2_X1 _10947_ ( .A1(_03773_ ), .A2(_03774_ ), .ZN(_03775_ ) );
AOI21_X1 _10948_ ( .A(_01940_ ), .B1(_03712_ ), .B2(_03713_ ), .ZN(_03776_ ) );
OAI21_X1 _10949_ ( .A(_01078_ ), .B1(_03775_ ), .B2(_03776_ ), .ZN(_03777_ ) );
AOI21_X1 _10950_ ( .A(_01076_ ), .B1(_03750_ ), .B2(_03777_ ), .ZN(_00167_ ) );
NOR2_X1 _10951_ ( .A1(_01996_ ), .A2(_03470_ ), .ZN(_03778_ ) );
OAI21_X2 _10952_ ( .A(_01054_ ), .B1(_03677_ ), .B2(_03778_ ), .ZN(_03779_ ) );
NOR2_X1 _10953_ ( .A1(\ar_data[16] ), .A2(_03492_ ), .ZN(_03780_ ) );
AOI22_X1 _10954_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03781_ ) );
NAND3_X1 _10955_ ( .A1(_03721_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03782_ ) );
NAND3_X1 _10956_ ( .A1(_03581_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03783_ ) );
NAND4_X1 _10957_ ( .A1(_03781_ ), .A2(_03621_ ), .A3(_03782_ ), .A4(_03783_ ), .ZN(_03784_ ) );
AOI22_X1 _10958_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03506_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03785_ ) );
NAND3_X1 _10959_ ( .A1(_03581_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03786_ ) );
NAND3_X1 _10960_ ( .A1(_03684_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03787_ ) );
NAND4_X1 _10961_ ( .A1(_03785_ ), .A2(_03505_ ), .A3(_03786_ ), .A4(_03787_ ), .ZN(_03788_ ) );
AND3_X1 _10962_ ( .A1(_03784_ ), .A2(_03788_ ), .A3(_01044_ ), .ZN(_03789_ ) );
AOI22_X1 _10963_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03790_ ) );
AOI21_X1 _10964_ ( .A(_03596_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03791_ ) );
NAND3_X1 _10965_ ( .A1(_03697_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03792_ ) );
NAND3_X1 _10966_ ( .A1(_03790_ ), .A2(_03791_ ), .A3(_03792_ ), .ZN(_03793_ ) );
NAND3_X1 _10967_ ( .A1(_03515_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03794_ ) );
NAND3_X1 _10968_ ( .A1(_03525_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03795_ ) );
NAND2_X1 _10969_ ( .A1(_03794_ ), .A2(_03795_ ), .ZN(_03796_ ) );
AOI21_X1 _10970_ ( .A(_03525_ ), .B1(\u_reg.rf[1][16] ), .B2(_03599_ ), .ZN(_03797_ ) );
OR3_X1 _10971_ ( .A1(_03796_ ), .A2(_03505_ ), .A3(_03797_ ), .ZN(_03798_ ) );
AND2_X1 _10972_ ( .A1(_03798_ ), .A2(_03705_ ), .ZN(_03799_ ) );
AOI21_X1 _10973_ ( .A(_03789_ ), .B1(_03793_ ), .B2(_03799_ ), .ZN(_03800_ ) );
OAI21_X1 _10974_ ( .A(_03681_ ), .B1(_03546_ ), .B2(_03800_ ), .ZN(_03801_ ) );
OAI21_X1 _10975_ ( .A(_03638_ ), .B1(_03780_ ), .B2(_03801_ ), .ZN(_03802_ ) );
NAND3_X1 _10976_ ( .A1(_01983_ ), .A2(_01989_ ), .A3(_03643_ ), .ZN(_03803_ ) );
AND3_X1 _10977_ ( .A1(_03802_ ), .A2(_03476_ ), .A3(_03803_ ), .ZN(_03804_ ) );
AOI21_X1 _10978_ ( .A(_01996_ ), .B1(_03712_ ), .B2(_03713_ ), .ZN(_03805_ ) );
OAI21_X1 _10979_ ( .A(_01078_ ), .B1(_03804_ ), .B2(_03805_ ), .ZN(_03806_ ) );
AOI21_X1 _10980_ ( .A(_01076_ ), .B1(_03779_ ), .B2(_03806_ ), .ZN(_00168_ ) );
BUF_X4 _10981_ ( .A(_01075_ ), .Z(_03807_ ) );
NOR2_X1 _10982_ ( .A1(_02037_ ), .A2(_03470_ ), .ZN(_03808_ ) );
OAI21_X2 _10983_ ( .A(_01054_ ), .B1(_03677_ ), .B2(_03808_ ), .ZN(_03809_ ) );
AOI22_X1 _10984_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03810_ ) );
NAND3_X1 _10985_ ( .A1(_03627_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03811_ ) );
NAND3_X1 _10986_ ( .A1(_03573_ ), .A2(_03574_ ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03812_ ) );
NAND4_X1 _10987_ ( .A1(_03810_ ), .A2(_03702_ ), .A3(_03811_ ), .A4(_03812_ ), .ZN(_03813_ ) );
AOI22_X1 _10988_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03814_ ) );
NAND3_X1 _10989_ ( .A1(_03609_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03815_ ) );
NAND3_X1 _10990_ ( .A1(_03609_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03816_ ) );
NAND4_X1 _10991_ ( .A1(_03814_ ), .A2(_03646_ ), .A3(_03815_ ), .A4(_03816_ ), .ZN(_03817_ ) );
NAND3_X1 _10992_ ( .A1(_03813_ ), .A2(_03817_ ), .A3(_03559_ ), .ZN(_03818_ ) );
AOI22_X1 _10993_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03506_ ), .B1(_03565_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03819_ ) );
NAND3_X1 _10994_ ( .A1(_03721_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03820_ ) );
NAND2_X1 _10995_ ( .A1(_03819_ ), .A2(_03820_ ), .ZN(_03821_ ) );
AOI211_X1 _10996_ ( .A(_03702_ ), .B(_03821_ ), .C1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03695_ ), .ZN(_03822_ ) );
NAND3_X1 _10997_ ( .A1(_03525_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03823_ ) );
INV_X1 _10998_ ( .A(_03565_ ), .ZN(_03824_ ) );
OAI21_X1 _10999_ ( .A(_03823_ ), .B1(_03824_ ), .B2(_02014_ ), .ZN(_03825_ ) );
AOI21_X1 _11000_ ( .A(_03606_ ), .B1(\u_reg.rf[1][15] ), .B2(_03599_ ), .ZN(_03826_ ) );
OR3_X1 _11001_ ( .A1(_03825_ ), .A2(_03505_ ), .A3(_03826_ ), .ZN(_03827_ ) );
NAND2_X1 _11002_ ( .A1(_03827_ ), .A2(_03705_ ), .ZN(_03828_ ) );
OAI21_X1 _11003_ ( .A(_03818_ ), .B1(_03822_ ), .B2(_03828_ ), .ZN(_03829_ ) );
AOI21_X1 _11004_ ( .A(_03482_ ), .B1(_03536_ ), .B2(_03829_ ), .ZN(_03830_ ) );
OAI21_X1 _11005_ ( .A(_03830_ ), .B1(\ar_data[15] ), .B2(_03492_ ), .ZN(_03831_ ) );
AOI21_X1 _11006_ ( .A(_03477_ ), .B1(_03831_ ), .B2(_03638_ ), .ZN(_03832_ ) );
NAND3_X1 _11007_ ( .A1(_02025_ ), .A2(_03589_ ), .A3(_02030_ ), .ZN(_03833_ ) );
AND2_X1 _11008_ ( .A1(_03832_ ), .A2(_03833_ ), .ZN(_03834_ ) );
AOI21_X1 _11009_ ( .A(_02037_ ), .B1(_03712_ ), .B2(_03713_ ), .ZN(_03835_ ) );
OAI21_X1 _11010_ ( .A(_01078_ ), .B1(_03834_ ), .B2(_03835_ ), .ZN(_03836_ ) );
AOI21_X1 _11011_ ( .A(_03807_ ), .B1(_03809_ ), .B2(_03836_ ), .ZN(_00169_ ) );
NOR2_X1 _11012_ ( .A1(_02090_ ), .A2(_03470_ ), .ZN(_03837_ ) );
OAI21_X2 _11013_ ( .A(_01054_ ), .B1(_03677_ ), .B2(_03837_ ), .ZN(_03838_ ) );
AOI22_X1 _11014_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03839_ ) );
NAND3_X1 _11015_ ( .A1(_03607_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03840_ ) );
NAND3_X1 _11016_ ( .A1(_03607_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03841_ ) );
NAND4_X1 _11017_ ( .A1(_03839_ ), .A2(_03702_ ), .A3(_03840_ ), .A4(_03841_ ), .ZN(_03842_ ) );
AOI21_X1 _11018_ ( .A(_03524_ ), .B1(_03531_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03843_ ) );
NAND3_X1 _11019_ ( .A1(_03627_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03844_ ) );
NAND3_X1 _11020_ ( .A1(_03609_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03845_ ) );
NAND3_X1 _11021_ ( .A1(_03603_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03846_ ) );
NAND4_X1 _11022_ ( .A1(_03843_ ), .A2(_03844_ ), .A3(_03845_ ), .A4(_03846_ ), .ZN(_03847_ ) );
NAND3_X1 _11023_ ( .A1(_03842_ ), .A2(_03559_ ), .A3(_03847_ ), .ZN(_03848_ ) );
AOI22_X1 _11024_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03849_ ) );
AOI22_X1 _11025_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03850_ ) );
NAND3_X1 _11026_ ( .A1(_03849_ ), .A2(_03850_ ), .A3(_03557_ ), .ZN(_03851_ ) );
NAND2_X1 _11027_ ( .A1(_03851_ ), .A2(_03614_ ), .ZN(_03852_ ) );
AND3_X1 _11028_ ( .A1(_03609_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03853_ ) );
AND3_X1 _11029_ ( .A1(_03721_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03854_ ) );
AOI21_X1 _11030_ ( .A(_03576_ ), .B1(\u_reg.rf[1][14] ), .B2(_03603_ ), .ZN(_03855_ ) );
NOR4_X1 _11031_ ( .A1(_03853_ ), .A2(_03854_ ), .A3(_03855_ ), .A4(_03570_ ), .ZN(_03856_ ) );
OAI21_X1 _11032_ ( .A(_03848_ ), .B1(_03852_ ), .B2(_03856_ ), .ZN(_03857_ ) );
AOI21_X1 _11033_ ( .A(_03482_ ), .B1(_03536_ ), .B2(_03857_ ), .ZN(_03858_ ) );
OAI21_X1 _11034_ ( .A(_03858_ ), .B1(\ar_data[14] ), .B2(_03492_ ), .ZN(_03859_ ) );
AOI21_X1 _11035_ ( .A(_03477_ ), .B1(_03859_ ), .B2(_03638_ ), .ZN(_03860_ ) );
NAND3_X1 _11036_ ( .A1(_02078_ ), .A2(_02084_ ), .A3(_03589_ ), .ZN(_03861_ ) );
AND2_X1 _11037_ ( .A1(_03860_ ), .A2(_03861_ ), .ZN(_03862_ ) );
NOR2_X1 _11038_ ( .A1(_02090_ ), .A2(_03746_ ), .ZN(_03863_ ) );
OAI21_X1 _11039_ ( .A(_01077_ ), .B1(_03862_ ), .B2(_03863_ ), .ZN(_03864_ ) );
AOI21_X1 _11040_ ( .A(_03807_ ), .B1(_03838_ ), .B2(_03864_ ), .ZN(_00170_ ) );
NOR2_X1 _11041_ ( .A1(_02136_ ), .A2(_03470_ ), .ZN(_03865_ ) );
OAI21_X2 _11042_ ( .A(_01054_ ), .B1(_03677_ ), .B2(_03865_ ), .ZN(_03866_ ) );
AOI22_X1 _11043_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03867_ ) );
NAND3_X1 _11044_ ( .A1(_03607_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03868_ ) );
NAND3_X1 _11045_ ( .A1(_03607_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03869_ ) );
NAND4_X1 _11046_ ( .A1(_03867_ ), .A2(_03702_ ), .A3(_03868_ ), .A4(_03869_ ), .ZN(_03870_ ) );
AOI21_X1 _11047_ ( .A(_03524_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03871_ ) );
NAND3_X1 _11048_ ( .A1(_03627_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03872_ ) );
NAND3_X1 _11049_ ( .A1(_03609_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03873_ ) );
NAND3_X1 _11050_ ( .A1(_03603_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03874_ ) );
NAND4_X1 _11051_ ( .A1(_03871_ ), .A2(_03872_ ), .A3(_03873_ ), .A4(_03874_ ), .ZN(_03875_ ) );
NAND3_X1 _11052_ ( .A1(_03870_ ), .A2(_03559_ ), .A3(_03875_ ), .ZN(_03876_ ) );
AOI22_X1 _11053_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03877_ ) );
AOI22_X1 _11054_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03878_ ) );
NAND3_X1 _11055_ ( .A1(_03877_ ), .A2(_03878_ ), .A3(_03632_ ), .ZN(_03879_ ) );
NAND2_X1 _11056_ ( .A1(_03879_ ), .A2(_03614_ ), .ZN(_03880_ ) );
AND3_X1 _11057_ ( .A1(_03576_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03881_ ) );
AND3_X1 _11058_ ( .A1(_03581_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03882_ ) );
AOI21_X1 _11059_ ( .A(_03721_ ), .B1(\u_reg.rf[1][13] ), .B2(_03603_ ), .ZN(_03883_ ) );
NOR4_X1 _11060_ ( .A1(_03881_ ), .A2(_03882_ ), .A3(_03883_ ), .A4(_03570_ ), .ZN(_03884_ ) );
OAI21_X1 _11061_ ( .A(_03876_ ), .B1(_03880_ ), .B2(_03884_ ), .ZN(_03885_ ) );
AOI21_X1 _11062_ ( .A(_03482_ ), .B1(_03536_ ), .B2(_03885_ ), .ZN(_03886_ ) );
OAI21_X1 _11063_ ( .A(_03886_ ), .B1(\ar_data[13] ), .B2(_03492_ ), .ZN(_03887_ ) );
AOI21_X1 _11064_ ( .A(_03477_ ), .B1(_03887_ ), .B2(_03638_ ), .ZN(_03888_ ) );
NAND3_X1 _11065_ ( .A1(_02124_ ), .A2(_02130_ ), .A3(_03589_ ), .ZN(_03889_ ) );
AND2_X1 _11066_ ( .A1(_03888_ ), .A2(_03889_ ), .ZN(_03890_ ) );
NOR2_X1 _11067_ ( .A1(_02136_ ), .A2(_03746_ ), .ZN(_03891_ ) );
OAI21_X1 _11068_ ( .A(_01077_ ), .B1(_03890_ ), .B2(_03891_ ), .ZN(_03892_ ) );
AOI21_X1 _11069_ ( .A(_03807_ ), .B1(_03866_ ), .B2(_03892_ ), .ZN(_00171_ ) );
NOR2_X1 _11070_ ( .A1(_02172_ ), .A2(_03470_ ), .ZN(_03893_ ) );
OAI21_X2 _11071_ ( .A(_01053_ ), .B1(_03677_ ), .B2(_03893_ ), .ZN(_03894_ ) );
NOR2_X1 _11072_ ( .A1(\ar_data[12] ), .A2(_03492_ ), .ZN(_03895_ ) );
AOI22_X1 _11073_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03506_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03896_ ) );
NAND3_X1 _11074_ ( .A1(_03688_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03897_ ) );
NAND3_X1 _11075_ ( .A1(_03650_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03898_ ) );
AND4_X1 _11076_ ( .A1(_03524_ ), .A2(_03896_ ), .A3(_03897_ ), .A4(_03898_ ), .ZN(_03899_ ) );
NAND3_X1 _11077_ ( .A1(_03515_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03900_ ) );
NAND2_X1 _11078_ ( .A1(_03900_ ), .A2(_03487_ ), .ZN(_03901_ ) );
NAND3_X1 _11079_ ( .A1(_03606_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03902_ ) );
NAND3_X1 _11080_ ( .A1(_03606_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03903_ ) );
NAND2_X1 _11081_ ( .A1(_03902_ ), .A2(_03903_ ), .ZN(_03904_ ) );
AOI211_X1 _11082_ ( .A(_03901_ ), .B(_03904_ ), .C1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03531_ ), .ZN(_03905_ ) );
NOR3_X1 _11083_ ( .A1(_03899_ ), .A2(_03905_ ), .A3(_03705_ ), .ZN(_03906_ ) );
AOI21_X1 _11084_ ( .A(_03596_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03907_ ) );
NAND3_X1 _11085_ ( .A1(_03697_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03908_ ) );
BUF_X4 _11086_ ( .A(_03603_ ), .Z(_03909_ ) );
NAND3_X1 _11087_ ( .A1(_03909_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03910_ ) );
NAND3_X1 _11088_ ( .A1(_03909_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03911_ ) );
NAND4_X1 _11089_ ( .A1(_03907_ ), .A2(_03908_ ), .A3(_03910_ ), .A4(_03911_ ), .ZN(_03912_ ) );
NAND3_X1 _11090_ ( .A1(_03519_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03913_ ) );
OAI21_X1 _11091_ ( .A(_03913_ ), .B1(_03824_ ), .B2(_02151_ ), .ZN(_03914_ ) );
OAI211_X1 _11092_ ( .A(fanout_net_22 ), .B(\u_reg.rf[1][12] ), .C1(_02689_ ), .C2(_00668_ ), .ZN(_03915_ ) );
AOI211_X1 _11093_ ( .A(_03570_ ), .B(_03914_ ), .C1(_03573_ ), .C2(_03915_ ), .ZN(_03916_ ) );
NOR2_X1 _11094_ ( .A1(_03916_ ), .A2(_03559_ ), .ZN(_03917_ ) );
AOI21_X1 _11095_ ( .A(_03906_ ), .B1(_03912_ ), .B2(_03917_ ), .ZN(_03918_ ) );
OAI21_X1 _11096_ ( .A(_03681_ ), .B1(_03546_ ), .B2(_03918_ ), .ZN(_03919_ ) );
OAI21_X1 _11097_ ( .A(_03638_ ), .B1(_03895_ ), .B2(_03919_ ), .ZN(_03920_ ) );
OR3_X1 _11098_ ( .A1(_02180_ ), .A2(_03540_ ), .A3(_02181_ ), .ZN(_03921_ ) );
AND3_X1 _11099_ ( .A1(_03920_ ), .A2(_03476_ ), .A3(_03921_ ), .ZN(_03922_ ) );
NOR2_X1 _11100_ ( .A1(_02172_ ), .A2(_02407_ ), .ZN(_03923_ ) );
OAI21_X1 _11101_ ( .A(_01077_ ), .B1(_03922_ ), .B2(_03923_ ), .ZN(_03924_ ) );
AOI21_X1 _11102_ ( .A(_03807_ ), .B1(_03894_ ), .B2(_03924_ ), .ZN(_00172_ ) );
AND3_X1 _11103_ ( .A1(_02209_ ), .A2(_03643_ ), .A3(_02215_ ), .ZN(_03925_ ) );
AOI21_X1 _11104_ ( .A(_03517_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03926_ ) );
NAND3_X1 _11105_ ( .A1(_03650_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03927_ ) );
NAND3_X1 _11106_ ( .A1(_03734_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03928_ ) );
NAND3_X1 _11107_ ( .A1(_03599_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03929_ ) );
AND4_X1 _11108_ ( .A1(_03926_ ), .A2(_03927_ ), .A3(_03928_ ), .A4(_03929_ ), .ZN(_03930_ ) );
AOI21_X1 _11109_ ( .A(_03632_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03931_ ) );
AND3_X1 _11110_ ( .A1(_03509_ ), .A2(_00875_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03932_ ) );
AOI221_X4 _11111_ ( .A(_03932_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03506_ ), .ZN(_03933_ ) );
AOI211_X1 _11112_ ( .A(_03705_ ), .B(_03930_ ), .C1(_03931_ ), .C2(_03933_ ), .ZN(_03934_ ) );
AOI22_X1 _11113_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03565_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03935_ ) );
BUF_X4 _11114_ ( .A(_03502_ ), .Z(_03936_ ) );
AOI22_X1 _11115_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03937_ ) );
AND3_X1 _11116_ ( .A1(_03935_ ), .A2(_03937_ ), .A3(_03570_ ), .ZN(_03938_ ) );
AND3_X1 _11117_ ( .A1(_03734_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03939_ ) );
AND3_X1 _11118_ ( .A1(_03606_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03940_ ) );
AOI21_X1 _11119_ ( .A(_03519_ ), .B1(\u_reg.rf[1][29] ), .B2(_03650_ ), .ZN(_03941_ ) );
NOR4_X1 _11120_ ( .A1(_03939_ ), .A2(_03940_ ), .A3(_03941_ ), .A4(_03505_ ), .ZN(_03942_ ) );
NOR3_X1 _11121_ ( .A1(_03938_ ), .A2(_03559_ ), .A3(_03942_ ), .ZN(_03943_ ) );
OR2_X1 _11122_ ( .A1(_03934_ ), .A2(_03943_ ), .ZN(_03944_ ) );
AOI21_X1 _11123_ ( .A(_03594_ ), .B1(_03537_ ), .B2(_03944_ ), .ZN(_03945_ ) );
AND2_X1 _11124_ ( .A1(_02187_ ), .A2(_02189_ ), .ZN(\ar_data[29] ) );
BUF_X4 _11125_ ( .A(_03536_ ), .Z(_03946_ ) );
OAI21_X1 _11126_ ( .A(_03945_ ), .B1(\ar_data[29] ), .B2(_03946_ ), .ZN(_03947_ ) );
AOI211_X1 _11127_ ( .A(_03478_ ), .B(_03925_ ), .C1(_03947_ ), .C2(_03541_ ), .ZN(_03948_ ) );
NOR2_X1 _11128_ ( .A1(_02219_ ), .A2(_03746_ ), .ZN(_03949_ ) );
OAI21_X1 _11129_ ( .A(_03592_ ), .B1(_03948_ ), .B2(_03949_ ), .ZN(_03950_ ) );
OAI21_X1 _11130_ ( .A(_03950_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00173_ ) );
BUF_X8 _11131_ ( .A(_03469_ ), .Z(_03951_ ) );
OAI211_X1 _11132_ ( .A(_01869_ ), .B(_02269_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_03952_ ) );
NAND3_X1 _11133_ ( .A1(_02256_ ), .A2(_02262_ ), .A3(_03589_ ), .ZN(_03953_ ) );
AND2_X1 _11134_ ( .A1(_02230_ ), .A2(_02232_ ), .ZN(\ar_data[11] ) );
OR2_X1 _11135_ ( .A1(\ar_data[11] ), .A2(_03536_ ), .ZN(_03954_ ) );
CLKBUF_X2 _11136_ ( .A(_03681_ ), .Z(_03955_ ) );
NAND3_X1 _11137_ ( .A1(_03515_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03956_ ) );
NAND3_X1 _11138_ ( .A1(_03497_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03957_ ) );
NAND3_X1 _11139_ ( .A1(_03494_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03958_ ) );
AND3_X1 _11140_ ( .A1(_03956_ ), .A2(_03957_ ), .A3(_03958_ ), .ZN(_03959_ ) );
AOI21_X1 _11141_ ( .A(_03487_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03960_ ) );
AOI21_X1 _11142_ ( .A(_03524_ ), .B1(_03531_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03961_ ) );
AND3_X1 _11143_ ( .A1(_03483_ ), .A2(_00875_ ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03962_ ) );
AOI221_X4 _11144_ ( .A(_03962_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_00996_ ), .ZN(_03963_ ) );
AOI221_X4 _11145_ ( .A(_03493_ ), .B1(_03959_ ), .B2(_03960_ ), .C1(_03961_ ), .C2(_03963_ ), .ZN(_03964_ ) );
AOI22_X1 _11146_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03965_ ) );
AOI22_X1 _11147_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03966_ ) );
NAND3_X1 _11148_ ( .A1(_03965_ ), .A2(_03966_ ), .A3(_03632_ ), .ZN(_03967_ ) );
OAI21_X1 _11149_ ( .A(_03573_ ), .B1(_03574_ ), .B2(_02246_ ), .ZN(_03968_ ) );
NAND3_X1 _11150_ ( .A1(_03607_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03969_ ) );
NAND3_X1 _11151_ ( .A1(_03607_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03970_ ) );
NAND4_X1 _11152_ ( .A1(_03968_ ), .A2(_03702_ ), .A3(_03969_ ), .A4(_03970_ ), .ZN(_03971_ ) );
AND3_X1 _11153_ ( .A1(_03967_ ), .A2(_03614_ ), .A3(_03971_ ), .ZN(_03972_ ) );
OAI21_X1 _11154_ ( .A(_03536_ ), .B1(_03964_ ), .B2(_03972_ ), .ZN(_03973_ ) );
AND3_X1 _11155_ ( .A1(_03954_ ), .A2(_03955_ ), .A3(_03973_ ), .ZN(_03974_ ) );
OAI211_X1 _11156_ ( .A(_03476_ ), .B(_03953_ ), .C1(_03974_ ), .C2(_03589_ ), .ZN(_03975_ ) );
OAI21_X1 _11157_ ( .A(_03975_ ), .B1(_03746_ ), .B2(_02268_ ), .ZN(_03976_ ) );
NAND2_X1 _11158_ ( .A1(_03976_ ), .A2(_00302_ ), .ZN(_03977_ ) );
NAND2_X1 _11159_ ( .A1(_03952_ ), .A2(_03977_ ), .ZN(_00174_ ) );
OAI211_X1 _11160_ ( .A(_01869_ ), .B(_02318_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_03978_ ) );
NOR2_X1 _11161_ ( .A1(\ar_data[10] ), .A2(_03537_ ), .ZN(_03979_ ) );
AOI22_X1 _11162_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03980_ ) );
NAND3_X1 _11163_ ( .A1(_03576_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03981_ ) );
NAND3_X1 _11164_ ( .A1(_03576_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03982_ ) );
NAND4_X1 _11165_ ( .A1(_03980_ ), .A2(_03621_ ), .A3(_03981_ ), .A4(_03982_ ), .ZN(_03983_ ) );
AOI22_X1 _11166_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03984_ ) );
NAND3_X1 _11167_ ( .A1(_03721_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03985_ ) );
NAND3_X1 _11168_ ( .A1(_03684_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03986_ ) );
NAND4_X1 _11169_ ( .A1(_03984_ ), .A2(_03570_ ), .A3(_03985_ ), .A4(_03986_ ), .ZN(_03987_ ) );
AND3_X1 _11170_ ( .A1(_03983_ ), .A2(_03987_ ), .A3(_01044_ ), .ZN(_03988_ ) );
NAND3_X1 _11171_ ( .A1(_03599_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03989_ ) );
NAND3_X1 _11172_ ( .A1(_03519_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03990_ ) );
NAND2_X1 _11173_ ( .A1(_03989_ ), .A2(_03990_ ), .ZN(_03991_ ) );
AOI21_X1 _11174_ ( .A(_03519_ ), .B1(\u_reg.rf[1][10] ), .B2(_03599_ ), .ZN(_03992_ ) );
OR3_X1 _11175_ ( .A1(_03991_ ), .A2(_03505_ ), .A3(_03992_ ), .ZN(_03993_ ) );
AND2_X1 _11176_ ( .A1(_03993_ ), .A2(_03614_ ), .ZN(_03994_ ) );
AOI22_X1 _11177_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03995_ ) );
AOI21_X1 _11178_ ( .A(_03596_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03996_ ) );
NAND3_X1 _11179_ ( .A1(_03697_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03997_ ) );
NAND3_X1 _11180_ ( .A1(_03995_ ), .A2(_03996_ ), .A3(_03997_ ), .ZN(_03998_ ) );
AOI21_X1 _11181_ ( .A(_03988_ ), .B1(_03994_ ), .B2(_03998_ ), .ZN(_03999_ ) );
OAI21_X1 _11182_ ( .A(_03681_ ), .B1(_03546_ ), .B2(_03999_ ), .ZN(_04000_ ) );
OAI21_X1 _11183_ ( .A(_03638_ ), .B1(_03979_ ), .B2(_04000_ ), .ZN(_04001_ ) );
NAND3_X1 _11184_ ( .A1(_02303_ ), .A2(_03589_ ), .A3(_02309_ ), .ZN(_04002_ ) );
AND3_X1 _11185_ ( .A1(_04001_ ), .A2(_03476_ ), .A3(_04002_ ), .ZN(_04003_ ) );
NOR2_X1 _11186_ ( .A1(_02317_ ), .A2(_03746_ ), .ZN(_04004_ ) );
OAI21_X1 _11187_ ( .A(_00302_ ), .B1(_04003_ ), .B2(_04004_ ), .ZN(_04005_ ) );
NAND2_X1 _11188_ ( .A1(_03978_ ), .A2(_04005_ ), .ZN(_00175_ ) );
NAND3_X1 _11189_ ( .A1(_01053_ ), .A2(_01060_ ), .A3(_02361_ ), .ZN(_04006_ ) );
NOR2_X1 _11190_ ( .A1(_03472_ ), .A2(_04006_ ), .ZN(_04007_ ) );
NAND3_X1 _11191_ ( .A1(_02350_ ), .A2(_03643_ ), .A3(_02355_ ), .ZN(_04008_ ) );
AND2_X1 _11192_ ( .A1(_02327_ ), .A2(_02329_ ), .ZN(\ar_data[9] ) );
OR2_X1 _11193_ ( .A1(\ar_data[9] ), .A2(_03491_ ), .ZN(_04009_ ) );
AOI21_X1 _11194_ ( .A(_03517_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04010_ ) );
NAND3_X1 _11195_ ( .A1(_03684_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04011_ ) );
NAND3_X1 _11196_ ( .A1(_03688_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04012_ ) );
NAND3_X1 _11197_ ( .A1(_03650_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04013_ ) );
AND4_X1 _11198_ ( .A1(_04010_ ), .A2(_04011_ ), .A3(_04012_ ), .A4(_04013_ ), .ZN(_04014_ ) );
AOI21_X1 _11199_ ( .A(_03557_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04015_ ) );
AND3_X1 _11200_ ( .A1(_03497_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04016_ ) );
AOI221_X4 _11201_ ( .A(_04016_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03506_ ), .ZN(_04017_ ) );
AOI211_X1 _11202_ ( .A(_03705_ ), .B(_04014_ ), .C1(_04015_ ), .C2(_04017_ ), .ZN(_04018_ ) );
AOI22_X1 _11203_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04019_ ) );
AOI22_X1 _11204_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04020_ ) );
AND3_X1 _11205_ ( .A1(_04019_ ), .A2(_04020_ ), .A3(_03646_ ), .ZN(_04021_ ) );
AND3_X1 _11206_ ( .A1(_03581_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04022_ ) );
AND3_X1 _11207_ ( .A1(_03734_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04023_ ) );
AOI21_X1 _11208_ ( .A(_03734_ ), .B1(\u_reg.rf[1][9] ), .B2(_03684_ ), .ZN(_04024_ ) );
NOR4_X1 _11209_ ( .A1(_04022_ ), .A2(_04023_ ), .A3(_04024_ ), .A4(_03505_ ), .ZN(_04025_ ) );
NOR3_X1 _11210_ ( .A1(_04021_ ), .A2(_03559_ ), .A3(_04025_ ), .ZN(_04026_ ) );
OAI21_X1 _11211_ ( .A(_03536_ ), .B1(_04018_ ), .B2(_04026_ ), .ZN(_04027_ ) );
AND3_X1 _11212_ ( .A1(_04009_ ), .A2(_03955_ ), .A3(_04027_ ), .ZN(_04028_ ) );
OAI211_X1 _11213_ ( .A(_03476_ ), .B(_04008_ ), .C1(_04028_ ), .C2(_03589_ ), .ZN(_04029_ ) );
NAND2_X1 _11214_ ( .A1(_01861_ ), .A2(_02361_ ), .ZN(_04030_ ) );
AOI21_X1 _11215_ ( .A(_01805_ ), .B1(_04029_ ), .B2(_04030_ ), .ZN(_04031_ ) );
OR2_X1 _11216_ ( .A1(_04007_ ), .A2(_04031_ ), .ZN(_00176_ ) );
OAI211_X1 _11217_ ( .A(_01869_ ), .B(_02405_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_04032_ ) );
AND3_X1 _11218_ ( .A1(_02395_ ), .A2(_03643_ ), .A3(_02401_ ), .ZN(_04033_ ) );
AND3_X1 _11219_ ( .A1(_03497_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04034_ ) );
AOI221_X4 _11220_ ( .A(_04034_ ), .B1(_03565_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03647_ ), .ZN(_04035_ ) );
NAND3_X1 _11221_ ( .A1(_03909_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04036_ ) );
NAND3_X1 _11222_ ( .A1(_04035_ ), .A2(_03622_ ), .A3(_04036_ ), .ZN(_04037_ ) );
AOI22_X1 _11223_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04038_ ) );
AOI22_X1 _11224_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04039_ ) );
NAND3_X1 _11225_ ( .A1(_04038_ ), .A2(_04039_ ), .A3(_03571_ ), .ZN(_04040_ ) );
NAND3_X1 _11226_ ( .A1(_04037_ ), .A2(_03662_ ), .A3(_04040_ ), .ZN(_04041_ ) );
AND3_X1 _11227_ ( .A1(_03734_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04042_ ) );
AND3_X1 _11228_ ( .A1(_03606_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04043_ ) );
AOI21_X1 _11229_ ( .A(_03734_ ), .B1(\u_reg.rf[1][8] ), .B2(_03650_ ), .ZN(_04044_ ) );
OR4_X1 _11230_ ( .A1(_03646_ ), .A2(_04042_ ), .A3(_04043_ ), .A4(_04044_ ), .ZN(_04045_ ) );
AOI22_X1 _11231_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04046_ ) );
AOI22_X1 _11232_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04047_ ) );
NAND3_X1 _11233_ ( .A1(_04046_ ), .A2(_04047_ ), .A3(_03571_ ), .ZN(_04048_ ) );
NAND2_X1 _11234_ ( .A1(_04045_ ), .A2(_04048_ ), .ZN(_04049_ ) );
OAI21_X1 _11235_ ( .A(_04041_ ), .B1(_03662_ ), .B2(_04049_ ), .ZN(_04050_ ) );
AOI21_X1 _11236_ ( .A(_03594_ ), .B1(_03946_ ), .B2(_04050_ ), .ZN(_04051_ ) );
OAI21_X1 _11237_ ( .A(_04051_ ), .B1(\ar_data[8] ), .B2(_03946_ ), .ZN(_04052_ ) );
AOI211_X1 _11238_ ( .A(_03545_ ), .B(_04033_ ), .C1(_04052_ ), .C2(_03639_ ), .ZN(_04053_ ) );
AOI221_X4 _11239_ ( .A(_00890_ ), .B1(_01470_ ), .B2(_02359_ ), .C1(_03713_ ), .C2(_03712_ ), .ZN(_04054_ ) );
OAI21_X1 _11240_ ( .A(_00302_ ), .B1(_04053_ ), .B2(_04054_ ), .ZN(_04055_ ) );
NAND2_X1 _11241_ ( .A1(_04032_ ), .A2(_04055_ ), .ZN(_00177_ ) );
OAI211_X1 _11242_ ( .A(_01869_ ), .B(_02408_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_04056_ ) );
NAND4_X1 _11243_ ( .A1(_01772_ ), .A2(_00822_ ), .A3(_00821_ ), .A4(_01773_ ), .ZN(_04057_ ) );
NAND3_X1 _11244_ ( .A1(_01424_ ), .A2(_01773_ ), .A3(_02441_ ), .ZN(_04058_ ) );
AND3_X1 _11245_ ( .A1(_04057_ ), .A2(_03643_ ), .A3(_04058_ ), .ZN(_04059_ ) );
AOI22_X1 _11246_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04060_ ) );
NAND3_X1 _11247_ ( .A1(_03577_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04061_ ) );
NAND3_X1 _11248_ ( .A1(_03577_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04062_ ) );
NAND4_X1 _11249_ ( .A1(_04060_ ), .A2(_03553_ ), .A3(_04061_ ), .A4(_04062_ ), .ZN(_04063_ ) );
AOI21_X1 _11250_ ( .A(_03621_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04064_ ) );
NAND3_X1 _11251_ ( .A1(_03577_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04065_ ) );
NAND3_X1 _11252_ ( .A1(_03651_ ), .A2(fanout_net_23 ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04066_ ) );
NAND3_X1 _11253_ ( .A1(_03651_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04067_ ) );
NAND4_X1 _11254_ ( .A1(_04064_ ), .A2(_04065_ ), .A3(_04066_ ), .A4(_04067_ ), .ZN(_04068_ ) );
NAND3_X1 _11255_ ( .A1(_04063_ ), .A2(_03662_ ), .A3(_04068_ ), .ZN(_04069_ ) );
AOI22_X1 _11256_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04070_ ) );
AOI22_X1 _11257_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04071_ ) );
NAND3_X1 _11258_ ( .A1(_04070_ ), .A2(_04071_ ), .A3(_03571_ ), .ZN(_04072_ ) );
NAND2_X1 _11259_ ( .A1(_04072_ ), .A2(_03561_ ), .ZN(_04073_ ) );
OAI21_X1 _11260_ ( .A(_03573_ ), .B1(_03574_ ), .B2(_02420_ ), .ZN(_04074_ ) );
NAND3_X1 _11261_ ( .A1(_03577_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04075_ ) );
NAND3_X1 _11262_ ( .A1(_03582_ ), .A2(fanout_net_22 ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04076_ ) );
AND4_X1 _11263_ ( .A1(_03553_ ), .A2(_04074_ ), .A3(_04075_ ), .A4(_04076_ ), .ZN(_04077_ ) );
OAI21_X1 _11264_ ( .A(_04069_ ), .B1(_04073_ ), .B2(_04077_ ), .ZN(_04078_ ) );
AOI21_X1 _11265_ ( .A(_03594_ ), .B1(_03537_ ), .B2(_04078_ ), .ZN(_04079_ ) );
BUF_X4 _11266_ ( .A(_03537_ ), .Z(_04080_ ) );
OAI21_X1 _11267_ ( .A(_04079_ ), .B1(\ar_data[7] ), .B2(_04080_ ), .ZN(_04081_ ) );
AOI211_X1 _11268_ ( .A(_03545_ ), .B(_04059_ ), .C1(_04081_ ), .C2(_03639_ ), .ZN(_04082_ ) );
AOI221_X4 _11269_ ( .A(_00707_ ), .B1(_01470_ ), .B2(_02359_ ), .C1(_03713_ ), .C2(_03712_ ), .ZN(_04083_ ) );
OAI21_X1 _11270_ ( .A(_00302_ ), .B1(_04082_ ), .B2(_04083_ ), .ZN(_04084_ ) );
NAND2_X1 _11271_ ( .A1(_04056_ ), .A2(_04084_ ), .ZN(_00178_ ) );
OAI211_X1 _11272_ ( .A(_01869_ ), .B(_02489_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_04085_ ) );
NOR3_X1 _11273_ ( .A1(_02483_ ), .A2(_03540_ ), .A3(_02484_ ), .ZN(_04086_ ) );
AOI22_X1 _11274_ ( .A1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04087_ ) );
NAND3_X1 _11275_ ( .A1(_03909_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04088_ ) );
NAND3_X1 _11276_ ( .A1(_03573_ ), .A2(_03574_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04089_ ) );
NAND4_X1 _11277_ ( .A1(_04087_ ), .A2(_03557_ ), .A3(_04088_ ), .A4(_04089_ ), .ZN(_04090_ ) );
AOI22_X1 _11278_ ( .A1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04091_ ) );
NAND3_X1 _11279_ ( .A1(_03577_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04092_ ) );
NAND3_X1 _11280_ ( .A1(_03577_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04093_ ) );
NAND4_X1 _11281_ ( .A1(_04091_ ), .A2(_03553_ ), .A3(_04092_ ), .A4(_04093_ ), .ZN(_04094_ ) );
NAND3_X1 _11282_ ( .A1(_04090_ ), .A2(_04094_ ), .A3(_03662_ ), .ZN(_04095_ ) );
AOI22_X1 _11283_ ( .A1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04096_ ) );
AOI21_X1 _11284_ ( .A(_03596_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04097_ ) );
NAND3_X1 _11285_ ( .A1(_03697_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04098_ ) );
AND3_X1 _11286_ ( .A1(_04096_ ), .A2(_04097_ ), .A3(_04098_ ), .ZN(_04099_ ) );
AND3_X1 _11287_ ( .A1(_03688_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04100_ ) );
AOI21_X1 _11288_ ( .A(_04100_ ), .B1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03566_ ), .ZN(_04101_ ) );
AND2_X1 _11289_ ( .A1(_03600_ ), .A2(\u_reg.rf[1][6] ), .ZN(_04102_ ) );
OAI211_X1 _11290_ ( .A(_04101_ ), .B(_03553_ ), .C1(_03624_ ), .C2(_04102_ ), .ZN(_04103_ ) );
NAND2_X1 _11291_ ( .A1(_04103_ ), .A2(_03561_ ), .ZN(_04104_ ) );
OAI21_X1 _11292_ ( .A(_04095_ ), .B1(_04099_ ), .B2(_04104_ ), .ZN(_04105_ ) );
AOI21_X1 _11293_ ( .A(_03594_ ), .B1(_03946_ ), .B2(_04105_ ), .ZN(_04106_ ) );
OAI21_X1 _11294_ ( .A(_04106_ ), .B1(\ar_data[6] ), .B2(_04080_ ), .ZN(_04107_ ) );
AOI211_X1 _11295_ ( .A(_03545_ ), .B(_04086_ ), .C1(_04107_ ), .C2(_03639_ ), .ZN(_04108_ ) );
AOI221_X4 _11296_ ( .A(_00880_ ), .B1(_01470_ ), .B2(_02359_ ), .C1(_01081_ ), .C2(_01465_ ), .ZN(_04109_ ) );
OAI21_X1 _11297_ ( .A(_00302_ ), .B1(_04108_ ), .B2(_04109_ ), .ZN(_04110_ ) );
NAND2_X1 _11298_ ( .A1(_04085_ ), .A2(_04110_ ), .ZN(_00179_ ) );
OAI211_X1 _11299_ ( .A(_01869_ ), .B(_02531_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_04111_ ) );
NOR3_X1 _11300_ ( .A1(_02525_ ), .A2(_03540_ ), .A3(_02526_ ), .ZN(_04112_ ) );
AND3_X1 _11301_ ( .A1(_03497_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04113_ ) );
AOI221_X4 _11302_ ( .A(_04113_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03936_ ), .ZN(_04114_ ) );
NAND3_X1 _11303_ ( .A1(_03909_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04115_ ) );
NAND3_X1 _11304_ ( .A1(_04114_ ), .A2(_03622_ ), .A3(_04115_ ), .ZN(_04116_ ) );
AOI22_X1 _11305_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04117_ ) );
NAND3_X1 _11306_ ( .A1(_03651_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04118_ ) );
NAND3_X1 _11307_ ( .A1(_03573_ ), .A2(_03574_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04119_ ) );
NAND4_X1 _11308_ ( .A1(_04117_ ), .A2(_03557_ ), .A3(_04118_ ), .A4(_04119_ ), .ZN(_04120_ ) );
NAND3_X1 _11309_ ( .A1(_04116_ ), .A2(_03662_ ), .A3(_04120_ ), .ZN(_04121_ ) );
AOI21_X1 _11310_ ( .A(_03702_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04122_ ) );
NAND3_X1 _11311_ ( .A1(_03577_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04123_ ) );
NAND3_X1 _11312_ ( .A1(_03909_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04124_ ) );
NAND3_X1 _11313_ ( .A1(_03651_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04125_ ) );
AND4_X1 _11314_ ( .A1(_04122_ ), .A2(_04123_ ), .A3(_04124_ ), .A4(_04125_ ), .ZN(_04126_ ) );
AND3_X1 _11315_ ( .A1(_03525_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04127_ ) );
AND3_X1 _11316_ ( .A1(_03515_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04128_ ) );
OR2_X1 _11317_ ( .A1(_04127_ ), .A2(_04128_ ), .ZN(_04129_ ) );
AOI21_X1 _11318_ ( .A(_03576_ ), .B1(\u_reg.rf[1][5] ), .B2(_03603_ ), .ZN(_04130_ ) );
OR3_X1 _11319_ ( .A1(_04129_ ), .A2(_03632_ ), .A3(_04130_ ), .ZN(_04131_ ) );
NAND2_X1 _11320_ ( .A1(_04131_ ), .A2(_03614_ ), .ZN(_04132_ ) );
OAI21_X1 _11321_ ( .A(_04121_ ), .B1(_04126_ ), .B2(_04132_ ), .ZN(_04133_ ) );
AOI21_X1 _11322_ ( .A(_03594_ ), .B1(_03537_ ), .B2(_04133_ ), .ZN(_04134_ ) );
OAI21_X1 _11323_ ( .A(_04134_ ), .B1(\ar_data[5] ), .B2(_04080_ ), .ZN(_04135_ ) );
AOI211_X1 _11324_ ( .A(_03545_ ), .B(_04112_ ), .C1(_04135_ ), .C2(_03639_ ), .ZN(_04136_ ) );
AOI221_X4 _11325_ ( .A(_00891_ ), .B1(_01470_ ), .B2(_02359_ ), .C1(_01081_ ), .C2(_01465_ ), .ZN(_04137_ ) );
OAI21_X1 _11326_ ( .A(_00302_ ), .B1(_04136_ ), .B2(_04137_ ), .ZN(_04138_ ) );
NAND2_X1 _11327_ ( .A1(_04111_ ), .A2(_04138_ ), .ZN(_00180_ ) );
OAI211_X1 _11328_ ( .A(_01869_ ), .B(_02583_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_04139_ ) );
AND3_X1 _11329_ ( .A1(_02567_ ), .A2(_03643_ ), .A3(_02572_ ), .ZN(_04140_ ) );
AND2_X1 _11330_ ( .A1(_02561_ ), .A2(_02563_ ), .ZN(\ar_data[4] ) );
OR2_X1 _11331_ ( .A1(\ar_data[4] ), .A2(_03492_ ), .ZN(_04141_ ) );
NAND3_X1 _11332_ ( .A1(_03752_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04142_ ) );
NAND3_X1 _11333_ ( .A1(_03627_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04143_ ) );
NAND3_X1 _11334_ ( .A1(_03627_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04144_ ) );
NAND3_X1 _11335_ ( .A1(_04142_ ), .A2(_04143_ ), .A3(_04144_ ), .ZN(_04145_ ) );
AOI211_X1 _11336_ ( .A(_03553_ ), .B(_04145_ ), .C1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03612_ ), .ZN(_04146_ ) );
AOI21_X1 _11337_ ( .A(_03571_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04147_ ) );
AND3_X1 _11338_ ( .A1(_03519_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04148_ ) );
AOI221_X4 _11339_ ( .A(_04148_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03507_ ), .ZN(_04149_ ) );
AOI211_X1 _11340_ ( .A(_03561_ ), .B(_04146_ ), .C1(_04147_ ), .C2(_04149_ ), .ZN(_04150_ ) );
AOI22_X1 _11341_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04151_ ) );
AOI22_X1 _11342_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04152_ ) );
AND3_X1 _11343_ ( .A1(_04151_ ), .A2(_04152_ ), .A3(_03571_ ), .ZN(_04153_ ) );
AND3_X1 _11344_ ( .A1(_03582_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04154_ ) );
AND3_X1 _11345_ ( .A1(_03752_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04155_ ) );
AOI21_X1 _11346_ ( .A(_03752_ ), .B1(\u_reg.rf[1][4] ), .B2(_03600_ ), .ZN(_04156_ ) );
NOR4_X1 _11347_ ( .A1(_04154_ ), .A2(_04155_ ), .A3(_04156_ ), .A4(_03557_ ), .ZN(_04157_ ) );
NOR3_X1 _11348_ ( .A1(_04153_ ), .A2(_03662_ ), .A3(_04157_ ), .ZN(_04158_ ) );
OAI21_X1 _11349_ ( .A(_03946_ ), .B1(_04150_ ), .B2(_04158_ ), .ZN(_04159_ ) );
NAND3_X1 _11350_ ( .A1(_04141_ ), .A2(_03955_ ), .A3(_04159_ ), .ZN(_04160_ ) );
AOI211_X1 _11351_ ( .A(_03545_ ), .B(_04140_ ), .C1(_04160_ ), .C2(_03639_ ), .ZN(_04161_ ) );
AOI22_X1 _11352_ ( .A1(_03713_ ), .A2(_03712_ ), .B1(_02581_ ), .B2(_02582_ ), .ZN(_04162_ ) );
OAI21_X1 _11353_ ( .A(_00302_ ), .B1(_04161_ ), .B2(_04162_ ), .ZN(_04163_ ) );
NAND2_X1 _11354_ ( .A1(_04139_ ), .A2(_04163_ ), .ZN(_00181_ ) );
OAI211_X1 _11355_ ( .A(_01869_ ), .B(_02639_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_04164_ ) );
AND4_X1 _11356_ ( .A1(_02628_ ), .A2(_01712_ ), .A3(_01425_ ), .A4(_01368_ ), .ZN(_04165_ ) );
NOR3_X1 _11357_ ( .A1(_02627_ ), .A2(_03540_ ), .A3(_04165_ ), .ZN(_04166_ ) );
AND3_X1 _11358_ ( .A1(_03497_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04167_ ) );
AOI221_X4 _11359_ ( .A(_04167_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03936_ ), .ZN(_04168_ ) );
NAND3_X1 _11360_ ( .A1(_03909_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04169_ ) );
NAND3_X1 _11361_ ( .A1(_04168_ ), .A2(_03622_ ), .A3(_04169_ ), .ZN(_04170_ ) );
AOI22_X1 _11362_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03507_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04171_ ) );
NAND3_X1 _11363_ ( .A1(_03577_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04172_ ) );
NAND3_X1 _11364_ ( .A1(_03651_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04173_ ) );
NAND4_X1 _11365_ ( .A1(_04171_ ), .A2(_03557_ ), .A3(_04172_ ), .A4(_04173_ ), .ZN(_04174_ ) );
NAND3_X1 _11366_ ( .A1(_04170_ ), .A2(_04174_ ), .A3(_03662_ ), .ZN(_04175_ ) );
AOI21_X1 _11367_ ( .A(_03702_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04176_ ) );
NAND3_X1 _11368_ ( .A1(_03697_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04177_ ) );
NAND3_X1 _11369_ ( .A1(_03909_ ), .A2(_01641_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04178_ ) );
NAND3_X1 _11370_ ( .A1(_03909_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04179_ ) );
AND4_X1 _11371_ ( .A1(_04176_ ), .A2(_04177_ ), .A3(_04178_ ), .A4(_04179_ ), .ZN(_04180_ ) );
AND3_X1 _11372_ ( .A1(_03688_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04181_ ) );
AOI21_X1 _11373_ ( .A(_04181_ ), .B1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03566_ ), .ZN(_04182_ ) );
AND2_X1 _11374_ ( .A1(_03600_ ), .A2(\u_reg.rf[1][3] ), .ZN(_04183_ ) );
OAI211_X1 _11375_ ( .A(_04182_ ), .B(_03553_ ), .C1(_03624_ ), .C2(_04183_ ), .ZN(_04184_ ) );
NAND2_X1 _11376_ ( .A1(_04184_ ), .A2(_03614_ ), .ZN(_04185_ ) );
OAI21_X1 _11377_ ( .A(_04175_ ), .B1(_04180_ ), .B2(_04185_ ), .ZN(_04186_ ) );
AOI21_X1 _11378_ ( .A(_03594_ ), .B1(_03946_ ), .B2(_04186_ ), .ZN(_04187_ ) );
OAI21_X1 _11379_ ( .A(_04187_ ), .B1(\ar_data[3] ), .B2(_04080_ ), .ZN(_04188_ ) );
AOI211_X1 _11380_ ( .A(_03545_ ), .B(_04166_ ), .C1(_04188_ ), .C2(_03639_ ), .ZN(_04189_ ) );
AOI21_X1 _11381_ ( .A(_02638_ ), .B1(_03712_ ), .B2(_03713_ ), .ZN(_04190_ ) );
OAI21_X1 _11382_ ( .A(_03592_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04191_ ) );
NAND2_X1 _11383_ ( .A1(_04164_ ), .A2(_04191_ ), .ZN(_00182_ ) );
AOI22_X1 _11384_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_00996_ ), .B1(_03502_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04192_ ) );
NAND3_X1 _11385_ ( .A1(_03509_ ), .A2(_00875_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04193_ ) );
NAND3_X1 _11386_ ( .A1(_00955_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04194_ ) );
AND4_X1 _11387_ ( .A1(_00972_ ), .A2(_04192_ ), .A3(_04193_ ), .A4(_04194_ ), .ZN(_04195_ ) );
NAND3_X1 _11388_ ( .A1(_00955_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04196_ ) );
NAND2_X1 _11389_ ( .A1(_04196_ ), .A2(_03487_ ), .ZN(_04197_ ) );
NAND3_X1 _11390_ ( .A1(_03483_ ), .A2(_00751_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04198_ ) );
NAND3_X1 _11391_ ( .A1(_03483_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04199_ ) );
NAND2_X1 _11392_ ( .A1(_04198_ ), .A2(_04199_ ), .ZN(_04200_ ) );
AOI211_X1 _11393_ ( .A(_04197_ ), .B(_04200_ ), .C1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03502_ ), .ZN(_04201_ ) );
OR3_X1 _11394_ ( .A1(_04195_ ), .A2(_04201_ ), .A3(_00971_ ), .ZN(_04202_ ) );
AOI22_X1 _11395_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_00996_ ), .B1(_03565_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04203_ ) );
AOI21_X1 _11396_ ( .A(_03517_ ), .B1(_03502_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04204_ ) );
NAND3_X1 _11397_ ( .A1(_03525_ ), .A2(_03498_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04205_ ) );
AND3_X1 _11398_ ( .A1(_04203_ ), .A2(_04204_ ), .A3(_04205_ ), .ZN(_04206_ ) );
AND3_X1 _11399_ ( .A1(_03509_ ), .A2(_00875_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04207_ ) );
AND3_X1 _11400_ ( .A1(_03483_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04208_ ) );
AOI21_X1 _11401_ ( .A(_03509_ ), .B1(\u_reg.rf[1][2] ), .B2(_03494_ ), .ZN(_04209_ ) );
OR3_X1 _11402_ ( .A1(_04207_ ), .A2(_04208_ ), .A3(_04209_ ), .ZN(_04210_ ) );
OAI21_X1 _11403_ ( .A(_03493_ ), .B1(_04210_ ), .B2(_03505_ ), .ZN(_04211_ ) );
OAI21_X1 _11404_ ( .A(_04202_ ), .B1(_04206_ ), .B2(_04211_ ), .ZN(_04212_ ) );
AOI21_X1 _11405_ ( .A(_03481_ ), .B1(_03491_ ), .B2(_04212_ ), .ZN(_04213_ ) );
OAI211_X1 _11406_ ( .A(_04213_ ), .B(_03539_ ), .C1(\ar_data[2] ), .C2(_03491_ ), .ZN(_04214_ ) );
OAI21_X1 _11407_ ( .A(_01418_ ), .B1(_02677_ ), .B2(_02683_ ), .ZN(_04215_ ) );
AOI21_X1 _11408_ ( .A(_03477_ ), .B1(_04214_ ), .B2(_04215_ ), .ZN(_04216_ ) );
AOI21_X1 _11409_ ( .A(_04216_ ), .B1(_01566_ ), .B2(_02693_ ), .ZN(_04217_ ) );
AND2_X1 _11410_ ( .A1(_03467_ ), .A2(_03468_ ), .ZN(_04218_ ) );
INV_X1 _11411_ ( .A(_04218_ ), .ZN(_04219_ ) );
OAI21_X1 _11412_ ( .A(_01452_ ), .B1(_04219_ ), .B2(_02693_ ), .ZN(_04220_ ) );
OR3_X1 _11413_ ( .A1(_02690_ ), .A2(_00747_ ), .A3(_02691_ ), .ZN(_04221_ ) );
AOI22_X1 _11414_ ( .A1(_01063_ ), .A2(_01066_ ), .B1(_03054_ ), .B2(_04221_ ), .ZN(_04222_ ) );
AOI221_X1 _11415_ ( .A(_00896_ ), .B1(_01077_ ), .B2(_04217_ ), .C1(_04220_ ), .C2(_04222_ ), .ZN(_00183_ ) );
NOR2_X1 _11416_ ( .A1(_02732_ ), .A2(_02407_ ), .ZN(_04223_ ) );
AOI21_X1 _11417_ ( .A(_03517_ ), .B1(_03502_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04224_ ) );
NAND3_X1 _11418_ ( .A1(_03509_ ), .A2(_00875_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04225_ ) );
NAND3_X1 _11419_ ( .A1(_03494_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04226_ ) );
NAND3_X1 _11420_ ( .A1(_03494_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04227_ ) );
AND3_X1 _11421_ ( .A1(_04225_ ), .A2(_04226_ ), .A3(_04227_ ), .ZN(_04228_ ) );
AND3_X1 _11422_ ( .A1(_03483_ ), .A2(_00751_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04229_ ) );
AOI221_X4 _11423_ ( .A(_04229_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_00996_ ), .ZN(_04230_ ) );
AOI21_X1 _11424_ ( .A(_03487_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04231_ ) );
AOI221_X4 _11425_ ( .A(_03493_ ), .B1(_04224_ ), .B2(_04228_ ), .C1(_04230_ ), .C2(_04231_ ), .ZN(_04232_ ) );
AOI22_X1 _11426_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04233_ ) );
AOI22_X1 _11427_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04234_ ) );
NAND3_X1 _11428_ ( .A1(_04233_ ), .A2(_04234_ ), .A3(_03570_ ), .ZN(_04235_ ) );
OAI21_X1 _11429_ ( .A(_00980_ ), .B1(_00981_ ), .B2(_02711_ ), .ZN(_04236_ ) );
NAND3_X1 _11430_ ( .A1(_03581_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04237_ ) );
NAND3_X1 _11431_ ( .A1(_03581_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04238_ ) );
NAND4_X1 _11432_ ( .A1(_04236_ ), .A2(_03621_ ), .A3(_04237_ ), .A4(_04238_ ), .ZN(_04239_ ) );
AND3_X1 _11433_ ( .A1(_04235_ ), .A2(_03493_ ), .A3(_04239_ ), .ZN(_04240_ ) );
OR2_X1 _11434_ ( .A1(_04232_ ), .A2(_04240_ ), .ZN(_04241_ ) );
AOI21_X1 _11435_ ( .A(_03482_ ), .B1(_03537_ ), .B2(_04241_ ), .ZN(_04242_ ) );
AND2_X1 _11436_ ( .A1(_02699_ ), .A2(_02701_ ), .ZN(\ar_data[28] ) );
OAI21_X1 _11437_ ( .A(_04242_ ), .B1(\ar_data[28] ), .B2(_03946_ ), .ZN(_04243_ ) );
AOI21_X1 _11438_ ( .A(_03545_ ), .B1(_04243_ ), .B2(_03541_ ), .ZN(_04244_ ) );
NAND3_X1 _11439_ ( .A1(_02722_ ), .A2(_02728_ ), .A3(_03589_ ), .ZN(_04245_ ) );
AOI21_X1 _11440_ ( .A(_04223_ ), .B1(_04244_ ), .B2(_04245_ ), .ZN(_04246_ ) );
OAI22_X1 _11441_ ( .A1(_03472_ ), .A2(_03474_ ), .B1(_01805_ ), .B2(_04246_ ), .ZN(_00184_ ) );
OAI211_X1 _11442_ ( .A(_01721_ ), .B(_02776_ ), .C1(_03951_ ), .C2(_03471_ ), .ZN(_04247_ ) );
NOR3_X1 _11443_ ( .A1(_02767_ ), .A2(_03540_ ), .A3(_02768_ ), .ZN(_04248_ ) );
AND3_X1 _11444_ ( .A1(_03721_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04249_ ) );
AOI21_X1 _11445_ ( .A(_04249_ ), .B1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03619_ ), .ZN(_04250_ ) );
AND2_X1 _11446_ ( .A1(_03651_ ), .A2(\u_reg.rf[1][1] ), .ZN(_04251_ ) );
OAI211_X1 _11447_ ( .A(_04250_ ), .B(_03622_ ), .C1(_03624_ ), .C2(_04251_ ), .ZN(_04252_ ) );
AOI22_X1 _11448_ ( .A1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03566_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04253_ ) );
AOI21_X1 _11449_ ( .A(_03596_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04254_ ) );
NAND3_X1 _11450_ ( .A1(_03697_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04255_ ) );
NAND3_X1 _11451_ ( .A1(_04253_ ), .A2(_04254_ ), .A3(_04255_ ), .ZN(_04256_ ) );
NAND3_X1 _11452_ ( .A1(_04252_ ), .A2(_03561_ ), .A3(_04256_ ), .ZN(_04257_ ) );
AOI22_X1 _11453_ ( .A1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04258_ ) );
NAND3_X1 _11454_ ( .A1(_03697_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04259_ ) );
NAND3_X1 _11455_ ( .A1(_03697_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04260_ ) );
NAND4_X1 _11456_ ( .A1(_04258_ ), .A2(_03622_ ), .A3(_04259_ ), .A4(_04260_ ), .ZN(_04261_ ) );
AOI22_X1 _11457_ ( .A1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03563_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04262_ ) );
NAND3_X1 _11458_ ( .A1(_03577_ ), .A2(_03698_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04263_ ) );
NAND3_X1 _11459_ ( .A1(_03909_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04264_ ) );
NAND4_X1 _11460_ ( .A1(_04262_ ), .A2(_03571_ ), .A3(_04263_ ), .A4(_04264_ ), .ZN(_04265_ ) );
NAND3_X1 _11461_ ( .A1(_04261_ ), .A2(_04265_ ), .A3(_03662_ ), .ZN(_04266_ ) );
NAND2_X1 _11462_ ( .A1(_04257_ ), .A2(_04266_ ), .ZN(_04267_ ) );
AOI21_X1 _11463_ ( .A(_03594_ ), .B1(_03537_ ), .B2(_04267_ ), .ZN(_04268_ ) );
OAI21_X1 _11464_ ( .A(_04268_ ), .B1(\ar_data[1] ), .B2(_03946_ ), .ZN(_04269_ ) );
AOI211_X1 _11465_ ( .A(_03545_ ), .B(_04248_ ), .C1(_04269_ ), .C2(_03639_ ), .ZN(_04270_ ) );
AOI22_X1 _11466_ ( .A1(_03713_ ), .A2(_03712_ ), .B1(_02774_ ), .B2(_02775_ ), .ZN(_04271_ ) );
OAI21_X1 _11467_ ( .A(_03592_ ), .B1(_04270_ ), .B2(_04271_ ), .ZN(_04272_ ) );
NAND2_X1 _11468_ ( .A1(_04247_ ), .A2(_04272_ ), .ZN(_00185_ ) );
AND3_X1 _11469_ ( .A1(_00720_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(_00687_ ), .ZN(_04273_ ) );
OAI211_X2 _11470_ ( .A(_01721_ ), .B(_02828_ ), .C1(_03951_ ), .C2(_04273_ ), .ZN(_04274_ ) );
NOR3_X1 _11471_ ( .A1(_02815_ ), .A2(_03540_ ), .A3(_02816_ ), .ZN(_04275_ ) );
AND2_X1 _11472_ ( .A1(_02805_ ), .A2(_02807_ ), .ZN(\ar_data[0] ) );
OR2_X1 _11473_ ( .A1(_03537_ ), .A2(\ar_data[0] ), .ZN(_04276_ ) );
NAND3_X1 _11474_ ( .A1(_03752_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04277_ ) );
NAND3_X1 _11475_ ( .A1(_03627_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04278_ ) );
NAND3_X1 _11476_ ( .A1(_03627_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04279_ ) );
NAND3_X1 _11477_ ( .A1(_04277_ ), .A2(_04278_ ), .A3(_04279_ ), .ZN(_04280_ ) );
AOI211_X1 _11478_ ( .A(_03596_ ), .B(_04280_ ), .C1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03612_ ), .ZN(_04281_ ) );
AOI21_X1 _11479_ ( .A(_03571_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04282_ ) );
AND3_X1 _11480_ ( .A1(_03599_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04283_ ) );
AOI221_X4 _11481_ ( .A(_04283_ ), .B1(_03522_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03507_ ), .ZN(_04284_ ) );
AOI211_X1 _11482_ ( .A(_03561_ ), .B(_04281_ ), .C1(_04282_ ), .C2(_04284_ ), .ZN(_04285_ ) );
AOI22_X1 _11483_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04286_ ) );
AOI22_X1 _11484_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03648_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04287_ ) );
AND3_X1 _11485_ ( .A1(_04286_ ), .A2(_04287_ ), .A3(_03571_ ), .ZN(_04288_ ) );
AND3_X1 _11486_ ( .A1(_03582_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04289_ ) );
AND3_X1 _11487_ ( .A1(_03752_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04290_ ) );
AOI21_X1 _11488_ ( .A(_03752_ ), .B1(\u_reg.rf[1][0] ), .B2(_03600_ ), .ZN(_04291_ ) );
NOR4_X1 _11489_ ( .A1(_04289_ ), .A2(_04290_ ), .A3(_04291_ ), .A4(_03557_ ), .ZN(_04292_ ) );
NOR3_X1 _11490_ ( .A1(_04288_ ), .A2(_03662_ ), .A3(_04292_ ), .ZN(_04293_ ) );
OAI21_X1 _11491_ ( .A(_03946_ ), .B1(_04285_ ), .B2(_04293_ ), .ZN(_04294_ ) );
NAND3_X1 _11492_ ( .A1(_04276_ ), .A2(_03955_ ), .A3(_04294_ ), .ZN(_04295_ ) );
AOI211_X1 _11493_ ( .A(_03545_ ), .B(_04275_ ), .C1(_04295_ ), .C2(_03639_ ), .ZN(_04296_ ) );
AOI21_X1 _11494_ ( .A(_02827_ ), .B1(_03713_ ), .B2(_03712_ ), .ZN(_04297_ ) );
OAI21_X1 _11495_ ( .A(_03592_ ), .B1(_04296_ ), .B2(_04297_ ), .ZN(_04298_ ) );
NAND2_X1 _11496_ ( .A1(_04274_ ), .A2(_04298_ ), .ZN(_00186_ ) );
AND3_X1 _11497_ ( .A1(_02858_ ), .A2(_03643_ ), .A3(_02864_ ), .ZN(_04299_ ) );
AOI22_X1 _11498_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03506_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04300_ ) );
NAND3_X1 _11499_ ( .A1(_03688_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04301_ ) );
NAND3_X1 _11500_ ( .A1(_03688_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04302_ ) );
AND4_X1 _11501_ ( .A1(_03621_ ), .A2(_04300_ ), .A3(_04301_ ), .A4(_04302_ ), .ZN(_04303_ ) );
NAND3_X1 _11502_ ( .A1(_03525_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04304_ ) );
NAND3_X1 _11503_ ( .A1(_03515_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04305_ ) );
NAND3_X1 _11504_ ( .A1(_03515_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04306_ ) );
NAND3_X1 _11505_ ( .A1(_04304_ ), .A2(_04305_ ), .A3(_04306_ ), .ZN(_04307_ ) );
AOI211_X1 _11506_ ( .A(_03524_ ), .B(_04307_ ), .C1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03531_ ), .ZN(_04308_ ) );
NOR3_X1 _11507_ ( .A1(_04303_ ), .A2(_04308_ ), .A3(_03705_ ), .ZN(_04309_ ) );
AND3_X1 _11508_ ( .A1(_03734_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04310_ ) );
AND3_X1 _11509_ ( .A1(_03519_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04311_ ) );
AOI21_X1 _11510_ ( .A(_03734_ ), .B1(\u_reg.rf[1][27] ), .B2(_03650_ ), .ZN(_04312_ ) );
OR4_X1 _11511_ ( .A1(_03632_ ), .A2(_04310_ ), .A3(_04311_ ), .A4(_04312_ ), .ZN(_04313_ ) );
AOI22_X1 _11512_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04314_ ) );
AOI22_X1 _11513_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04315_ ) );
NAND3_X1 _11514_ ( .A1(_04314_ ), .A2(_04315_ ), .A3(_03632_ ), .ZN(_04316_ ) );
AND2_X1 _11515_ ( .A1(_04316_ ), .A2(_03705_ ), .ZN(_04317_ ) );
AOI21_X1 _11516_ ( .A(_04309_ ), .B1(_04313_ ), .B2(_04317_ ), .ZN(_04318_ ) );
MUX2_X1 _11517_ ( .A(_04318_ ), .B(\ar_data[27] ), .S(_03546_ ), .Z(_04319_ ) );
NAND2_X1 _11518_ ( .A1(_04319_ ), .A2(_03955_ ), .ZN(_04320_ ) );
AOI211_X1 _11519_ ( .A(_03478_ ), .B(_04299_ ), .C1(_04320_ ), .C2(_03541_ ), .ZN(_04321_ ) );
NOR2_X1 _11520_ ( .A1(_02868_ ), .A2(_03746_ ), .ZN(_04322_ ) );
OAI21_X1 _11521_ ( .A(_03592_ ), .B1(_04321_ ), .B2(_04322_ ), .ZN(_04323_ ) );
OAI21_X1 _11522_ ( .A(_04323_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00187_ ) );
AND3_X1 _11523_ ( .A1(_02897_ ), .A2(_01418_ ), .A3(_02902_ ), .ZN(_04324_ ) );
AOI21_X1 _11524_ ( .A(_03594_ ), .B1(_02894_ ), .B2(_03548_ ), .ZN(_04325_ ) );
AOI22_X1 _11525_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03507_ ), .B1(_03531_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04326_ ) );
NAND3_X1 _11526_ ( .A1(_03752_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04327_ ) );
NAND3_X1 _11527_ ( .A1(_03600_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04328_ ) );
AND4_X1 _11528_ ( .A1(_03596_ ), .A2(_04326_ ), .A3(_04327_ ), .A4(_04328_ ), .ZN(_04329_ ) );
NAND3_X1 _11529_ ( .A1(_03603_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04330_ ) );
NAND2_X1 _11530_ ( .A1(_04330_ ), .A2(_03570_ ), .ZN(_04331_ ) );
NAND3_X1 _11531_ ( .A1(_03607_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04332_ ) );
NAND3_X1 _11532_ ( .A1(_03609_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04333_ ) );
NAND2_X1 _11533_ ( .A1(_04332_ ), .A2(_04333_ ), .ZN(_04334_ ) );
AOI211_X1 _11534_ ( .A(_04331_ ), .B(_04334_ ), .C1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03612_ ), .ZN(_04335_ ) );
NOR3_X1 _11535_ ( .A1(_04329_ ), .A2(_04335_ ), .A3(_03614_ ), .ZN(_04336_ ) );
NAND3_X1 _11536_ ( .A1(_03576_ ), .A2(_03629_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04337_ ) );
OAI21_X1 _11537_ ( .A(_04337_ ), .B1(_03824_ ), .B2(_02884_ ), .ZN(_04338_ ) );
AOI21_X1 _11538_ ( .A(_03609_ ), .B1(\u_reg.rf[1][26] ), .B2(_03600_ ), .ZN(_04339_ ) );
OR3_X1 _11539_ ( .A1(_04338_ ), .A2(_03632_ ), .A3(_04339_ ), .ZN(_04340_ ) );
AND2_X1 _11540_ ( .A1(_04340_ ), .A2(_03561_ ), .ZN(_04341_ ) );
AOI22_X1 _11541_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04342_ ) );
AOI21_X1 _11542_ ( .A(_03622_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04343_ ) );
NAND3_X1 _11543_ ( .A1(_03624_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04344_ ) );
NAND3_X1 _11544_ ( .A1(_04342_ ), .A2(_04343_ ), .A3(_04344_ ), .ZN(_04345_ ) );
AOI21_X1 _11545_ ( .A(_04336_ ), .B1(_04341_ ), .B2(_04345_ ), .ZN(_04346_ ) );
OAI21_X1 _11546_ ( .A(_04325_ ), .B1(_03548_ ), .B2(_04346_ ), .ZN(_04347_ ) );
AOI211_X1 _11547_ ( .A(_03478_ ), .B(_04324_ ), .C1(_04347_ ), .C2(_03541_ ), .ZN(_04348_ ) );
NOR2_X1 _11548_ ( .A1(_02906_ ), .A2(_03746_ ), .ZN(_04349_ ) );
OAI21_X1 _11549_ ( .A(_03592_ ), .B1(_04348_ ), .B2(_04349_ ), .ZN(_04350_ ) );
OAI21_X1 _11550_ ( .A(_04350_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00188_ ) );
AND3_X1 _11551_ ( .A1(_02935_ ), .A2(_01418_ ), .A3(_02940_ ), .ZN(_04351_ ) );
AOI21_X1 _11552_ ( .A(_03482_ ), .B1(_02932_ ), .B2(_03548_ ), .ZN(_04352_ ) );
AOI22_X1 _11553_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03568_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04353_ ) );
NAND3_X1 _11554_ ( .A1(_03651_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04354_ ) );
NAND3_X1 _11555_ ( .A1(_03573_ ), .A2(_03574_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04355_ ) );
NAND4_X1 _11556_ ( .A1(_04353_ ), .A2(_03557_ ), .A3(_04354_ ), .A4(_04355_ ), .ZN(_04356_ ) );
AOI22_X1 _11557_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03507_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04357_ ) );
NAND3_X1 _11558_ ( .A1(_03582_ ), .A2(_03579_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04358_ ) );
NAND3_X1 _11559_ ( .A1(_03582_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04359_ ) );
NAND4_X1 _11560_ ( .A1(_04357_ ), .A2(_03553_ ), .A3(_04358_ ), .A4(_04359_ ), .ZN(_04360_ ) );
AND3_X1 _11561_ ( .A1(_04356_ ), .A2(_04360_ ), .A3(_03559_ ), .ZN(_04361_ ) );
AOI22_X1 _11562_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04362_ ) );
AOI21_X1 _11563_ ( .A(_03622_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04363_ ) );
NAND3_X1 _11564_ ( .A1(_03624_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04364_ ) );
NAND3_X1 _11565_ ( .A1(_04362_ ), .A2(_04363_ ), .A3(_04364_ ), .ZN(_04365_ ) );
AND3_X1 _11566_ ( .A1(_03581_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04366_ ) );
AOI21_X1 _11567_ ( .A(_04366_ ), .B1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03619_ ), .ZN(_04367_ ) );
AND2_X1 _11568_ ( .A1(_03600_ ), .A2(\u_reg.rf[1][25] ), .ZN(_04368_ ) );
OAI211_X1 _11569_ ( .A(_04367_ ), .B(_03622_ ), .C1(_03624_ ), .C2(_04368_ ), .ZN(_04369_ ) );
AND2_X1 _11570_ ( .A1(_04369_ ), .A2(_03561_ ), .ZN(_04370_ ) );
AOI21_X1 _11571_ ( .A(_04361_ ), .B1(_04365_ ), .B2(_04370_ ), .ZN(_04371_ ) );
OAI21_X1 _11572_ ( .A(_04352_ ), .B1(_03548_ ), .B2(_04371_ ), .ZN(_04372_ ) );
AOI211_X1 _11573_ ( .A(_03478_ ), .B(_04351_ ), .C1(_04372_ ), .C2(_03541_ ), .ZN(_04373_ ) );
NOR2_X1 _11574_ ( .A1(_02944_ ), .A2(_03746_ ), .ZN(_04374_ ) );
OAI21_X1 _11575_ ( .A(_03592_ ), .B1(_04373_ ), .B2(_04374_ ), .ZN(_04375_ ) );
OAI21_X1 _11576_ ( .A(_04375_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00189_ ) );
NOR3_X1 _11577_ ( .A1(_02977_ ), .A2(_03540_ ), .A3(_02978_ ), .ZN(_04376_ ) );
AOI21_X1 _11578_ ( .A(_03517_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04377_ ) );
NAND3_X1 _11579_ ( .A1(_03734_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04378_ ) );
NAND3_X1 _11580_ ( .A1(_03599_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04379_ ) );
NAND3_X1 _11581_ ( .A1(_03599_ ), .A2(_01639_ ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04380_ ) );
AND4_X1 _11582_ ( .A1(_04377_ ), .A2(_04378_ ), .A3(_04379_ ), .A4(_04380_ ), .ZN(_04381_ ) );
AOI21_X1 _11583_ ( .A(_03632_ ), .B1(_03695_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04382_ ) );
AND3_X1 _11584_ ( .A1(_03509_ ), .A2(_00875_ ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04383_ ) );
AOI221_X4 _11585_ ( .A(_04383_ ), .B1(_03512_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03506_ ), .ZN(_04384_ ) );
AOI211_X1 _11586_ ( .A(_03705_ ), .B(_04381_ ), .C1(_04382_ ), .C2(_04384_ ), .ZN(_04385_ ) );
AOI22_X1 _11587_ ( .A1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04386_ ) );
AOI22_X1 _11588_ ( .A1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04387_ ) );
NAND3_X1 _11589_ ( .A1(_04386_ ), .A2(_04387_ ), .A3(_03646_ ), .ZN(_04388_ ) );
OAI21_X1 _11590_ ( .A(_00980_ ), .B1(_00981_ ), .B2(_02961_ ), .ZN(_04389_ ) );
NAND3_X1 _11591_ ( .A1(_03721_ ), .A2(_03722_ ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04390_ ) );
NAND3_X1 _11592_ ( .A1(_03721_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04391_ ) );
NAND4_X1 _11593_ ( .A1(_04389_ ), .A2(_03621_ ), .A3(_04390_ ), .A4(_04391_ ), .ZN(_04392_ ) );
AND3_X1 _11594_ ( .A1(_04388_ ), .A2(_03493_ ), .A3(_04392_ ), .ZN(_04393_ ) );
OR2_X1 _11595_ ( .A1(_04385_ ), .A2(_04393_ ), .ZN(_04394_ ) );
AOI21_X1 _11596_ ( .A(_03482_ ), .B1(_03537_ ), .B2(_04394_ ), .ZN(_04395_ ) );
AND2_X1 _11597_ ( .A1(_02949_ ), .A2(_02951_ ), .ZN(\ar_data[24] ) );
OAI21_X1 _11598_ ( .A(_04395_ ), .B1(\ar_data[24] ), .B2(_03946_ ), .ZN(_04396_ ) );
AOI211_X1 _11599_ ( .A(_03478_ ), .B(_04376_ ), .C1(_04396_ ), .C2(_03541_ ), .ZN(_04397_ ) );
NOR2_X1 _11600_ ( .A1(_02983_ ), .A2(_03746_ ), .ZN(_04398_ ) );
OAI21_X1 _11601_ ( .A(_03592_ ), .B1(_04397_ ), .B2(_04398_ ), .ZN(_04399_ ) );
OAI21_X1 _11602_ ( .A(_04399_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00190_ ) );
AND3_X1 _11603_ ( .A1(_03013_ ), .A2(_01418_ ), .A3(_03018_ ), .ZN(_04400_ ) );
AOI21_X1 _11604_ ( .A(_03482_ ), .B1(_03010_ ), .B2(_03546_ ), .ZN(_04401_ ) );
AOI22_X1 _11605_ ( .A1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03522_ ), .B1(_03618_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04402_ ) );
NAND3_X1 _11606_ ( .A1(_03600_ ), .A2(_03652_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04403_ ) );
NAND3_X1 _11607_ ( .A1(_03573_ ), .A2(_03574_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04404_ ) );
NAND4_X1 _11608_ ( .A1(_04402_ ), .A2(_03632_ ), .A3(_04403_ ), .A4(_04404_ ), .ZN(_04405_ ) );
AOI22_X1 _11609_ ( .A1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03616_ ), .B1(_03503_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04406_ ) );
NAND3_X1 _11610_ ( .A1(_03752_ ), .A2(_00877_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04407_ ) );
NAND3_X1 _11611_ ( .A1(_03752_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04408_ ) );
NAND4_X1 _11612_ ( .A1(_04406_ ), .A2(_03702_ ), .A3(_04407_ ), .A4(_04408_ ), .ZN(_04409_ ) );
AND3_X1 _11613_ ( .A1(_04405_ ), .A2(_04409_ ), .A3(_03559_ ), .ZN(_04410_ ) );
AOI22_X1 _11614_ ( .A1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03617_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04411_ ) );
AOI21_X1 _11615_ ( .A(_03553_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04412_ ) );
NAND3_X1 _11616_ ( .A1(_03624_ ), .A2(_00878_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04413_ ) );
NAND3_X1 _11617_ ( .A1(_04411_ ), .A2(_04412_ ), .A3(_04413_ ), .ZN(_04414_ ) );
AND3_X1 _11618_ ( .A1(_03606_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04415_ ) );
AOI21_X1 _11619_ ( .A(_04415_ ), .B1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03618_ ), .ZN(_04416_ ) );
AOI211_X1 _11620_ ( .A(_03722_ ), .B(_02994_ ), .C1(_00917_ ), .C2(_00693_ ), .ZN(_04417_ ) );
OAI211_X1 _11621_ ( .A(_04416_ ), .B(_03596_ ), .C1(_03697_ ), .C2(_04417_ ), .ZN(_04418_ ) );
AND2_X1 _11622_ ( .A1(_04418_ ), .A2(_03614_ ), .ZN(_04419_ ) );
AOI21_X1 _11623_ ( .A(_04410_ ), .B1(_04414_ ), .B2(_04419_ ), .ZN(_04420_ ) );
OAI21_X1 _11624_ ( .A(_04401_ ), .B1(_03548_ ), .B2(_04420_ ), .ZN(_04421_ ) );
AOI211_X1 _11625_ ( .A(_03478_ ), .B(_04400_ ), .C1(_04421_ ), .C2(_03541_ ), .ZN(_04422_ ) );
AOI21_X1 _11626_ ( .A(_04422_ ), .B1(_01861_ ), .B2(_03022_ ), .ZN(_04423_ ) );
OAI22_X1 _11627_ ( .A1(_03472_ ), .A2(_03474_ ), .B1(_01805_ ), .B2(_04423_ ), .ZN(_00191_ ) );
AND3_X1 _11628_ ( .A1(_03061_ ), .A2(_01418_ ), .A3(_03062_ ), .ZN(_04424_ ) );
AOI21_X1 _11629_ ( .A(_03536_ ), .B1(_03045_ ), .B2(_03047_ ), .ZN(_04425_ ) );
AOI22_X1 _11630_ ( .A1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03506_ ), .B1(_03530_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04426_ ) );
NAND3_X1 _11631_ ( .A1(_03581_ ), .A2(_03689_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04427_ ) );
NAND3_X1 _11632_ ( .A1(_03688_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04428_ ) );
NAND4_X1 _11633_ ( .A1(_04426_ ), .A2(_03621_ ), .A3(_04427_ ), .A4(_04428_ ), .ZN(_04429_ ) );
AOI21_X1 _11634_ ( .A(_03517_ ), .B1(_03936_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04430_ ) );
NAND3_X1 _11635_ ( .A1(_03684_ ), .A2(_01640_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04431_ ) );
NAND3_X1 _11636_ ( .A1(_03688_ ), .A2(_03578_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04432_ ) );
NAND3_X1 _11637_ ( .A1(_03650_ ), .A2(\u_idu.imm_auipc_lui[21] ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04433_ ) );
NAND4_X1 _11638_ ( .A1(_04430_ ), .A2(_04431_ ), .A3(_04432_ ), .A4(_04433_ ), .ZN(_04434_ ) );
AND3_X1 _11639_ ( .A1(_04429_ ), .A2(_01044_ ), .A3(_04434_ ), .ZN(_04435_ ) );
AND3_X1 _11640_ ( .A1(_03519_ ), .A2(_00876_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04436_ ) );
AND3_X1 _11641_ ( .A1(_03606_ ), .A2(\u_idu.imm_auipc_lui[20] ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04437_ ) );
AOI21_X1 _11642_ ( .A(_03519_ ), .B1(\u_reg.rf[1][22] ), .B2(_03650_ ), .ZN(_04438_ ) );
OR4_X1 _11643_ ( .A1(_03646_ ), .A2(_04436_ ), .A3(_04437_ ), .A4(_04438_ ), .ZN(_04439_ ) );
AOI22_X1 _11644_ ( .A1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03521_ ), .B1(_03549_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04440_ ) );
AOI22_X1 _11645_ ( .A1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03562_ ), .B1(_03647_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04441_ ) );
NAND3_X1 _11646_ ( .A1(_04440_ ), .A2(_04441_ ), .A3(_03646_ ), .ZN(_04442_ ) );
AND2_X1 _11647_ ( .A1(_04442_ ), .A2(_03493_ ), .ZN(_04443_ ) );
AOI21_X1 _11648_ ( .A(_04435_ ), .B1(_04439_ ), .B2(_04443_ ), .ZN(_04444_ ) );
OAI21_X1 _11649_ ( .A(_03681_ ), .B1(_03546_ ), .B2(_04444_ ), .ZN(_04445_ ) );
OR2_X1 _11650_ ( .A1(_04425_ ), .A2(_04445_ ), .ZN(_04446_ ) );
AOI211_X1 _11651_ ( .A(_03478_ ), .B(_04424_ ), .C1(_04446_ ), .C2(_03541_ ), .ZN(_04447_ ) );
AND2_X1 _11652_ ( .A1(_03051_ ), .A2(_01861_ ), .ZN(_04448_ ) );
OAI21_X1 _11653_ ( .A(_01804_ ), .B1(_04447_ ), .B2(_04448_ ), .ZN(_04449_ ) );
OAI21_X1 _11654_ ( .A(_04449_ ), .B1(_03473_ ), .B2(_03475_ ), .ZN(_00192_ ) );
AND3_X1 _11655_ ( .A1(_00865_ ), .A2(_00866_ ), .A3(_00946_ ), .ZN(_00193_ ) );
BUF_X4 _11656_ ( .A(_00856_ ), .Z(_04450_ ) );
NOR3_X1 _11657_ ( .A1(flush_$_OR__Y_B ), .A2(_00933_ ), .A3(_04450_ ), .ZN(_00194_ ) );
NOR3_X1 _11658_ ( .A1(flush_$_OR__Y_B ), .A2(_00937_ ), .A3(_04450_ ), .ZN(_00195_ ) );
NOR3_X1 _11659_ ( .A1(flush_$_OR__Y_B ), .A2(_00941_ ), .A3(_04450_ ), .ZN(_00196_ ) );
AOI21_X1 _11660_ ( .A(_03807_ ), .B1(_01422_ ), .B2(_01445_ ), .ZN(_00197_ ) );
AOI21_X1 _11661_ ( .A(_03807_ ), .B1(_01536_ ), .B2(_01552_ ), .ZN(_00198_ ) );
BUF_X4 _11662_ ( .A(_00896_ ), .Z(_04451_ ) );
BUF_X4 _11663_ ( .A(_04451_ ), .Z(_04452_ ) );
NOR2_X1 _11664_ ( .A1(_01635_ ), .A2(_04452_ ), .ZN(_00199_ ) );
AOI21_X1 _11665_ ( .A(_03807_ ), .B1(_01696_ ), .B2(_01714_ ), .ZN(_00200_ ) );
AOI21_X1 _11666_ ( .A(_03807_ ), .B1(_01774_ ), .B2(_01789_ ), .ZN(_00201_ ) );
AOI21_X1 _11667_ ( .A(_03807_ ), .B1(_01871_ ), .B2(_01878_ ), .ZN(_00202_ ) );
AOI21_X1 _11668_ ( .A(_03807_ ), .B1(_01932_ ), .B2(_01933_ ), .ZN(_00203_ ) );
BUF_X4 _11669_ ( .A(_01075_ ), .Z(_04453_ ) );
AOI21_X1 _11670_ ( .A(_04453_ ), .B1(_01983_ ), .B2(_01989_ ), .ZN(_00204_ ) );
AOI21_X1 _11671_ ( .A(_04453_ ), .B1(_02025_ ), .B2(_02030_ ), .ZN(_00205_ ) );
AOI21_X1 _11672_ ( .A(_04453_ ), .B1(_02078_ ), .B2(_02084_ ), .ZN(_00206_ ) );
AOI21_X1 _11673_ ( .A(_04453_ ), .B1(_02124_ ), .B2(_02130_ ), .ZN(_00207_ ) );
NOR2_X1 _11674_ ( .A1(_02182_ ), .A2(_04452_ ), .ZN(_00208_ ) );
AOI21_X1 _11675_ ( .A(_04453_ ), .B1(_02209_ ), .B2(_02215_ ), .ZN(_00209_ ) );
AOI21_X1 _11676_ ( .A(_04453_ ), .B1(_02256_ ), .B2(_02262_ ), .ZN(_00210_ ) );
AOI21_X1 _11677_ ( .A(_04453_ ), .B1(_02303_ ), .B2(_02309_ ), .ZN(_00211_ ) );
AOI21_X1 _11678_ ( .A(_04453_ ), .B1(_02350_ ), .B2(_02355_ ), .ZN(_00212_ ) );
AOI21_X1 _11679_ ( .A(_04453_ ), .B1(_02395_ ), .B2(_02401_ ), .ZN(_00213_ ) );
AOI21_X1 _11680_ ( .A(_04453_ ), .B1(_04057_ ), .B2(_04058_ ), .ZN(_00214_ ) );
NOR2_X1 _11681_ ( .A1(_02485_ ), .A2(_04452_ ), .ZN(_00215_ ) );
NOR2_X1 _11682_ ( .A1(_02527_ ), .A2(_04452_ ), .ZN(_00216_ ) );
BUF_X4 _11683_ ( .A(_01075_ ), .Z(_04454_ ) );
AOI21_X1 _11684_ ( .A(_04454_ ), .B1(_02567_ ), .B2(_02572_ ), .ZN(_00217_ ) );
NOR2_X1 _11685_ ( .A1(_02631_ ), .A2(_04452_ ), .ZN(_00218_ ) );
NOR2_X1 _11686_ ( .A1(_02684_ ), .A2(_04452_ ), .ZN(_00219_ ) );
AOI21_X1 _11687_ ( .A(_04454_ ), .B1(_02722_ ), .B2(_02728_ ), .ZN(_00220_ ) );
NOR2_X1 _11688_ ( .A1(_02769_ ), .A2(_04452_ ), .ZN(_00221_ ) );
NOR2_X1 _11689_ ( .A1(_02817_ ), .A2(_04452_ ), .ZN(_00222_ ) );
AOI21_X1 _11690_ ( .A(_04454_ ), .B1(_02858_ ), .B2(_02864_ ), .ZN(_00223_ ) );
AOI21_X1 _11691_ ( .A(_04454_ ), .B1(_02897_ ), .B2(_02902_ ), .ZN(_00224_ ) );
AOI21_X1 _11692_ ( .A(_04454_ ), .B1(_02935_ ), .B2(_02940_ ), .ZN(_00225_ ) );
NOR2_X1 _11693_ ( .A1(_02979_ ), .A2(_04452_ ), .ZN(_00226_ ) );
AOI21_X1 _11694_ ( .A(_04454_ ), .B1(_03013_ ), .B2(_03018_ ), .ZN(_00227_ ) );
AOI21_X1 _11695_ ( .A(_04454_ ), .B1(_03061_ ), .B2(_03062_ ), .ZN(_00228_ ) );
BUF_X4 _11696_ ( .A(_00856_ ), .Z(_04455_ ) );
BUF_X4 _11697_ ( .A(_00874_ ), .Z(_04456_ ) );
NOR3_X1 _11698_ ( .A1(_01105_ ), .A2(_04455_ ), .A3(_04456_ ), .ZN(_00232_ ) );
NOR3_X1 _11699_ ( .A1(flush_$_OR__Y_B ), .A2(_04455_ ), .A3(_01098_ ), .ZN(_00233_ ) );
AND4_X1 _11700_ ( .A1(_00674_ ), .A2(_00669_ ), .A3(_01097_ ), .A4(_03470_ ), .ZN(_04457_ ) );
AOI21_X1 _11701_ ( .A(_04454_ ), .B1(_04457_ ), .B2(_00739_ ), .ZN(_00234_ ) );
AND3_X1 _11702_ ( .A1(_00865_ ), .A2(\de_pc[31] ), .A3(_00866_ ), .ZN(_00235_ ) );
AND3_X1 _11703_ ( .A1(_00865_ ), .A2(\de_pc[30] ), .A3(_00866_ ), .ZN(_00236_ ) );
AND3_X1 _11704_ ( .A1(_00865_ ), .A2(\de_pc[21] ), .A3(_00866_ ), .ZN(_00237_ ) );
AND3_X1 _11705_ ( .A1(_00865_ ), .A2(\de_pc[20] ), .A3(_00866_ ), .ZN(_00238_ ) );
NOR4_X1 _11706_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_01792_ ), .ZN(_00239_ ) );
NOR4_X1 _11707_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_00860_ ), .A4(_01859_ ), .ZN(_00240_ ) );
BUF_X4 _11708_ ( .A(_00859_ ), .Z(_04458_ ) );
NOR4_X1 _11709_ ( .A1(_00861_ ), .A2(fanout_net_1 ), .A3(_04458_ ), .A4(_01935_ ), .ZN(_00241_ ) );
BUF_X4 _11710_ ( .A(_00856_ ), .Z(_04459_ ) );
NOR4_X1 _11711_ ( .A1(_04459_ ), .A2(fanout_net_1 ), .A3(_04458_ ), .A4(_01991_ ), .ZN(_00242_ ) );
NOR4_X1 _11712_ ( .A1(_04459_ ), .A2(fanout_net_1 ), .A3(_04458_ ), .A4(_02032_ ), .ZN(_00243_ ) );
NOR4_X1 _11713_ ( .A1(_04459_ ), .A2(fanout_net_1 ), .A3(_04458_ ), .A4(_02086_ ), .ZN(_00244_ ) );
NOR4_X1 _11714_ ( .A1(_04459_ ), .A2(fanout_net_1 ), .A3(_04458_ ), .A4(_02132_ ), .ZN(_00245_ ) );
NOR4_X1 _11715_ ( .A1(_04459_ ), .A2(fanout_net_2 ), .A3(_04458_ ), .A4(_02170_ ), .ZN(_00246_ ) );
CLKBUF_X2 _11716_ ( .A(_00637_ ), .Z(_04460_ ) );
AND3_X1 _11717_ ( .A1(_00865_ ), .A2(\de_pc[29] ), .A3(_04460_ ), .ZN(_00247_ ) );
AND3_X1 _11718_ ( .A1(_00865_ ), .A2(\de_pc[11] ), .A3(_04460_ ), .ZN(_00248_ ) );
NOR4_X1 _11719_ ( .A1(_04459_ ), .A2(fanout_net_2 ), .A3(_04458_ ), .A4(_02311_ ), .ZN(_00249_ ) );
AND3_X1 _11720_ ( .A1(_00865_ ), .A2(\de_pc[9] ), .A3(_04460_ ), .ZN(_00250_ ) );
AND3_X1 _11721_ ( .A1(_00865_ ), .A2(\de_pc[8] ), .A3(_04460_ ), .ZN(_00251_ ) );
NOR4_X1 _11722_ ( .A1(_04459_ ), .A2(fanout_net_2 ), .A3(_04458_ ), .A4(_02410_ ), .ZN(_00252_ ) );
CLKBUF_X2 _11723_ ( .A(_00864_ ), .Z(_04461_ ) );
AND3_X1 _11724_ ( .A1(_04461_ ), .A2(\de_pc[6] ), .A3(_04460_ ), .ZN(_00253_ ) );
AND3_X1 _11725_ ( .A1(_04461_ ), .A2(\de_pc[5] ), .A3(_04460_ ), .ZN(_00254_ ) );
NOR4_X1 _11726_ ( .A1(_04459_ ), .A2(fanout_net_2 ), .A3(_04458_ ), .A4(_02574_ ), .ZN(_00255_ ) );
NOR4_X1 _11727_ ( .A1(_04459_ ), .A2(fanout_net_2 ), .A3(_04458_ ), .A4(_02632_ ), .ZN(_00256_ ) );
BUF_X4 _11728_ ( .A(_00859_ ), .Z(_04462_ ) );
NOR4_X1 _11729_ ( .A1(_04459_ ), .A2(fanout_net_2 ), .A3(_04462_ ), .A4(_02685_ ), .ZN(_00257_ ) );
AND3_X1 _11730_ ( .A1(_04461_ ), .A2(\de_pc[28] ), .A3(_04460_ ), .ZN(_00258_ ) );
BUF_X4 _11731_ ( .A(_00856_ ), .Z(_04463_ ) );
NOR4_X1 _11732_ ( .A1(_04463_ ), .A2(fanout_net_2 ), .A3(_04462_ ), .A4(_02770_ ), .ZN(_00259_ ) );
NOR4_X1 _11733_ ( .A1(_04463_ ), .A2(fanout_net_2 ), .A3(_04462_ ), .A4(_02818_ ), .ZN(_00260_ ) );
AND3_X1 _11734_ ( .A1(_04461_ ), .A2(\de_pc[27] ), .A3(_04460_ ), .ZN(_00261_ ) );
AND3_X1 _11735_ ( .A1(_04461_ ), .A2(\de_pc[26] ), .A3(_04460_ ), .ZN(_00262_ ) );
AND3_X1 _11736_ ( .A1(_04461_ ), .A2(\de_pc[25] ), .A3(_04460_ ), .ZN(_00263_ ) );
CLKBUF_X2 _11737_ ( .A(_00637_ ), .Z(_04464_ ) );
AND3_X1 _11738_ ( .A1(_04461_ ), .A2(\de_pc[24] ), .A3(_04464_ ), .ZN(_00264_ ) );
AND3_X1 _11739_ ( .A1(_04461_ ), .A2(\de_pc[23] ), .A3(_04464_ ), .ZN(_00265_ ) );
NOR4_X1 _11740_ ( .A1(_04463_ ), .A2(fanout_net_2 ), .A3(_04462_ ), .A4(_03065_ ), .ZN(_00266_ ) );
NAND4_X1 _11741_ ( .A1(_00710_ ), .A2(_00868_ ), .A3(_00711_ ), .A4(_00713_ ), .ZN(_04465_ ) );
NOR4_X1 _11742_ ( .A1(flush_$_OR__Y_B ), .A2(_04450_ ), .A3(_00701_ ), .A4(_04465_ ), .ZN(_00267_ ) );
NOR4_X1 _11743_ ( .A1(_04463_ ), .A2(fanout_net_2 ), .A3(_04462_ ), .A4(_04465_ ), .ZN(_00268_ ) );
NOR2_X1 _11744_ ( .A1(_03538_ ), .A2(_04452_ ), .ZN(_00269_ ) );
BUF_X4 _11745_ ( .A(_04451_ ), .Z(_04466_ ) );
NOR2_X1 _11746_ ( .A1(_03587_ ), .A2(_04466_ ), .ZN(_00270_ ) );
NOR2_X1 _11747_ ( .A1(_03637_ ), .A2(_04466_ ), .ZN(_00271_ ) );
NOR2_X1 _11748_ ( .A1(_03673_ ), .A2(_04466_ ), .ZN(_00272_ ) );
BUF_X4 _11749_ ( .A(_01075_ ), .Z(_04467_ ) );
NOR3_X1 _11750_ ( .A1(_03680_ ), .A2(_04467_ ), .A3(_03708_ ), .ZN(_00273_ ) );
NOR3_X1 _11751_ ( .A1(_03718_ ), .A2(_04467_ ), .A3(_03742_ ), .ZN(_00274_ ) );
NOR2_X1 _11752_ ( .A1(_03772_ ), .A2(_04466_ ), .ZN(_00275_ ) );
NOR3_X1 _11753_ ( .A1(_03780_ ), .A2(_04467_ ), .A3(_03801_ ), .ZN(_00276_ ) );
NOR2_X1 _11754_ ( .A1(_03831_ ), .A2(_04466_ ), .ZN(_00277_ ) );
NOR2_X1 _11755_ ( .A1(_03859_ ), .A2(_04466_ ), .ZN(_00278_ ) );
NOR2_X1 _11756_ ( .A1(_03887_ ), .A2(_04466_ ), .ZN(_00279_ ) );
NOR3_X1 _11757_ ( .A1(_03895_ ), .A2(_01076_ ), .A3(_03919_ ), .ZN(_00280_ ) );
NOR2_X1 _11758_ ( .A1(_03947_ ), .A2(_04466_ ), .ZN(_00281_ ) );
AND4_X1 _11759_ ( .A1(_01061_ ), .A2(_03954_ ), .A3(_03955_ ), .A4(_03973_ ), .ZN(_00282_ ) );
NOR3_X1 _11760_ ( .A1(_03979_ ), .A2(_01076_ ), .A3(_04000_ ), .ZN(_00283_ ) );
AND4_X1 _11761_ ( .A1(_01061_ ), .A2(_04009_ ), .A3(_03955_ ), .A4(_04027_ ), .ZN(_00284_ ) );
NOR2_X1 _11762_ ( .A1(_04052_ ), .A2(_04466_ ), .ZN(_00285_ ) );
BUF_X2 _11763_ ( .A(_01060_ ), .Z(_04468_ ) );
OAI211_X1 _11764_ ( .A(_04468_ ), .B(_04079_ ), .C1(\ar_data[7] ), .C2(_04080_ ), .ZN(_04469_ ) );
INV_X1 _11765_ ( .A(_04469_ ), .ZN(_00286_ ) );
OAI211_X1 _11766_ ( .A(_04106_ ), .B(_04468_ ), .C1(\ar_data[6] ), .C2(_04080_ ), .ZN(_04470_ ) );
INV_X1 _11767_ ( .A(_04470_ ), .ZN(_00287_ ) );
OAI211_X1 _11768_ ( .A(_04468_ ), .B(_04134_ ), .C1(\ar_data[5] ), .C2(_04080_ ), .ZN(_04471_ ) );
INV_X1 _11769_ ( .A(_04471_ ), .ZN(_00288_ ) );
AND4_X1 _11770_ ( .A1(_01061_ ), .A2(_04141_ ), .A3(_03955_ ), .A4(_04159_ ), .ZN(_00289_ ) );
OAI211_X1 _11771_ ( .A(_04187_ ), .B(_04468_ ), .C1(\ar_data[3] ), .C2(_04080_ ), .ZN(_04472_ ) );
INV_X1 _11772_ ( .A(_04472_ ), .ZN(_00290_ ) );
OAI211_X1 _11773_ ( .A(_04213_ ), .B(_04468_ ), .C1(\ar_data[2] ), .C2(_04080_ ), .ZN(_04473_ ) );
INV_X1 _11774_ ( .A(_04473_ ), .ZN(_00291_ ) );
NOR2_X1 _11775_ ( .A1(_04243_ ), .A2(_04466_ ), .ZN(_00292_ ) );
OAI211_X1 _11776_ ( .A(_04268_ ), .B(_04468_ ), .C1(\ar_data[1] ), .C2(_04080_ ), .ZN(_04474_ ) );
INV_X1 _11777_ ( .A(_04474_ ), .ZN(_00293_ ) );
AND4_X1 _11778_ ( .A1(_01061_ ), .A2(_04276_ ), .A3(_03955_ ), .A4(_04294_ ), .ZN(_00294_ ) );
AND3_X1 _11779_ ( .A1(_04319_ ), .A2(_04468_ ), .A3(_03955_ ), .ZN(_00295_ ) );
BUF_X4 _11780_ ( .A(_04451_ ), .Z(_04475_ ) );
NOR2_X1 _11781_ ( .A1(_04347_ ), .A2(_04475_ ), .ZN(_00296_ ) );
NOR2_X1 _11782_ ( .A1(_04372_ ), .A2(_04475_ ), .ZN(_00297_ ) );
NOR2_X1 _11783_ ( .A1(_04396_ ), .A2(_04475_ ), .ZN(_00298_ ) );
NOR2_X1 _11784_ ( .A1(_04421_ ), .A2(_04475_ ), .ZN(_00299_ ) );
NOR3_X1 _11785_ ( .A1(_04425_ ), .A2(_01076_ ), .A3(_04445_ ), .ZN(_00300_ ) );
NOR2_X1 _11786_ ( .A1(_01025_ ), .A2(exu_valid ), .ZN(\u_exu.exe_end_$_ANDNOT__B_Y ) );
INV_X1 _11787_ ( .A(\u_exu.exe_end_$_ANDNOT__B_Y ), .ZN(_04476_ ) );
NOR4_X1 _11788_ ( .A1(_04463_ ), .A2(fanout_net_2 ), .A3(_04462_ ), .A4(_04476_ ), .ZN(_00301_ ) );
AND2_X1 _11789_ ( .A1(_03078_ ), .A2(fanout_net_20 ), .ZN(_04477_ ) );
BUF_X4 _11790_ ( .A(_04477_ ), .Z(_04478_ ) );
AOI21_X1 _11791_ ( .A(_03362_ ), .B1(_03358_ ), .B2(_03364_ ), .ZN(_04479_ ) );
OAI21_X1 _11792_ ( .A(_04478_ ), .B1(_03365_ ), .B2(_04479_ ), .ZN(_04480_ ) );
AND2_X1 _11793_ ( .A1(_03079_ ), .A2(\u_exu.alu_p1[5] ), .ZN(_04481_ ) );
BUF_X2 _11794_ ( .A(_03413_ ), .Z(_04482_ ) );
BUF_X2 _11795_ ( .A(_04482_ ), .Z(_04483_ ) );
AND2_X1 _11796_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[4] ), .ZN(_04484_ ) );
OR3_X1 _11797_ ( .A1(_04481_ ), .A2(_04483_ ), .A3(_04484_ ), .ZN(_04485_ ) );
AND2_X1 _11798_ ( .A1(_03080_ ), .A2(\u_exu.alu_p1[7] ), .ZN(_04486_ ) );
AND2_X1 _11799_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[6] ), .ZN(_04487_ ) );
OR3_X1 _11800_ ( .A1(_04486_ ), .A2(fanout_net_15 ), .A3(_04487_ ), .ZN(_04488_ ) );
BUF_X4 _11801_ ( .A(_03455_ ), .Z(_04489_ ) );
BUF_X2 _11802_ ( .A(_04489_ ), .Z(_04490_ ) );
NAND3_X1 _11803_ ( .A1(_04485_ ), .A2(_04488_ ), .A3(_04490_ ), .ZN(_04491_ ) );
AOI21_X1 _11804_ ( .A(_03463_ ), .B1(_03080_ ), .B2(\u_exu.alu_p1[1] ), .ZN(_04492_ ) );
AND2_X1 _11805_ ( .A1(_03079_ ), .A2(\u_exu.alu_p1[3] ), .ZN(_04493_ ) );
AND2_X1 _11806_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[2] ), .ZN(_04494_ ) );
NOR2_X1 _11807_ ( .A1(_04493_ ), .A2(_04494_ ), .ZN(_04495_ ) );
BUF_X2 _11808_ ( .A(_04482_ ), .Z(_04496_ ) );
MUX2_X1 _11809_ ( .A(_04492_ ), .B(_04495_ ), .S(_04496_ ), .Z(_04497_ ) );
BUF_X2 _11810_ ( .A(_03457_ ), .Z(_04498_ ) );
OAI211_X1 _11811_ ( .A(fanout_net_19 ), .B(_04491_ ), .C1(_04497_ ), .C2(_04498_ ), .ZN(_04499_ ) );
AND2_X2 _11812_ ( .A1(_03378_ ), .A2(\u_exu.alu_p2[4] ), .ZN(_04500_ ) );
BUF_X2 _11813_ ( .A(_04500_ ), .Z(_04501_ ) );
BUF_X4 _11814_ ( .A(_04496_ ), .Z(_04502_ ) );
AND2_X1 _11815_ ( .A1(_03079_ ), .A2(\u_exu.alu_p1[11] ), .ZN(_04503_ ) );
AND2_X1 _11816_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[10] ), .ZN(_04504_ ) );
OAI21_X1 _11817_ ( .A(_04502_ ), .B1(_04503_ ), .B2(_04504_ ), .ZN(_04505_ ) );
AND2_X1 _11818_ ( .A1(_03079_ ), .A2(\u_exu.alu_p1[9] ), .ZN(_04506_ ) );
AND2_X1 _11819_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[8] ), .ZN(_04507_ ) );
OAI21_X1 _11820_ ( .A(fanout_net_15 ), .B1(_04506_ ), .B2(_04507_ ), .ZN(_04508_ ) );
NAND2_X1 _11821_ ( .A1(_04505_ ), .A2(_04508_ ), .ZN(_04509_ ) );
NAND2_X1 _11822_ ( .A1(_04509_ ), .A2(fanout_net_17 ), .ZN(_04510_ ) );
AND2_X1 _11823_ ( .A1(_03080_ ), .A2(\u_exu.alu_p1[15] ), .ZN(_04511_ ) );
AND2_X1 _11824_ ( .A1(\u_exu.alu_p1[14] ), .A2(fanout_net_14 ), .ZN(_04512_ ) );
OR3_X1 _11825_ ( .A1(_04511_ ), .A2(fanout_net_15 ), .A3(_04512_ ), .ZN(_04513_ ) );
NOR2_X1 _11826_ ( .A1(_03192_ ), .A2(fanout_net_14 ), .ZN(_04514_ ) );
AND2_X1 _11827_ ( .A1(\u_exu.alu_p1[12] ), .A2(fanout_net_14 ), .ZN(_04515_ ) );
OR3_X1 _11828_ ( .A1(_04514_ ), .A2(_04515_ ), .A3(_04483_ ), .ZN(_04516_ ) );
NAND3_X1 _11829_ ( .A1(_04513_ ), .A2(_04498_ ), .A3(_04516_ ), .ZN(_04517_ ) );
BUF_X4 _11830_ ( .A(_03453_ ), .Z(_04518_ ) );
BUF_X4 _11831_ ( .A(_04518_ ), .Z(_04519_ ) );
BUF_X2 _11832_ ( .A(_04519_ ), .Z(_04520_ ) );
NAND3_X1 _11833_ ( .A1(_04510_ ), .A2(_04517_ ), .A3(_04520_ ), .ZN(_04521_ ) );
NAND3_X1 _11834_ ( .A1(_04499_ ), .A2(_04501_ ), .A3(_04521_ ), .ZN(_04522_ ) );
BUF_X4 _11835_ ( .A(_03454_ ), .Z(_04523_ ) );
BUF_X2 _11836_ ( .A(_04523_ ), .Z(_04524_ ) );
NOR2_X1 _11837_ ( .A1(_03347_ ), .A2(fanout_net_14 ), .ZN(_04525_ ) );
AND2_X1 _11838_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[28] ), .ZN(_04526_ ) );
NOR2_X1 _11839_ ( .A1(_04525_ ), .A2(_04526_ ), .ZN(_04527_ ) );
BUF_X2 _11840_ ( .A(_04483_ ), .Z(_04528_ ) );
NOR2_X1 _11841_ ( .A1(_04527_ ), .A2(_04528_ ), .ZN(_04529_ ) );
NOR2_X1 _11842_ ( .A1(_03361_ ), .A2(fanout_net_14 ), .ZN(_04530_ ) );
AND2_X1 _11843_ ( .A1(_04530_ ), .A2(_04502_ ), .ZN(_04531_ ) );
AND3_X1 _11844_ ( .A1(_04528_ ), .A2(\u_exu.alu_p1[30] ), .A3(fanout_net_14 ), .ZN(_04532_ ) );
NOR4_X1 _11845_ ( .A1(_04529_ ), .A2(fanout_net_17 ), .A3(_04531_ ), .A4(_04532_ ), .ZN(_04533_ ) );
AND2_X1 _11846_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[26] ), .ZN(_04534_ ) );
INV_X1 _11847_ ( .A(_04534_ ), .ZN(_04535_ ) );
OAI211_X1 _11848_ ( .A(_04535_ ), .B(_04528_ ), .C1(fanout_net_14 ), .C2(_03317_ ), .ZN(_04536_ ) );
NOR2_X1 _11849_ ( .A1(_03329_ ), .A2(fanout_net_14 ), .ZN(_04537_ ) );
INV_X1 _11850_ ( .A(_04537_ ), .ZN(_04538_ ) );
AND2_X1 _11851_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[24] ), .ZN(_04539_ ) );
INV_X1 _11852_ ( .A(_04539_ ), .ZN(_04540_ ) );
NAND3_X1 _11853_ ( .A1(_04538_ ), .A2(fanout_net_15 ), .A3(_04540_ ), .ZN(_04541_ ) );
AOI21_X1 _11854_ ( .A(_04498_ ), .B1(_04536_ ), .B2(_04541_ ), .ZN(_04542_ ) );
OAI21_X1 _11855_ ( .A(_04524_ ), .B1(_04533_ ), .B2(_04542_ ), .ZN(_04543_ ) );
AND2_X1 _11856_ ( .A1(_03080_ ), .A2(\u_exu.alu_p1[19] ), .ZN(_04544_ ) );
AND2_X1 _11857_ ( .A1(\u_exu.alu_p1[18] ), .A2(fanout_net_14 ), .ZN(_04545_ ) );
OAI21_X1 _11858_ ( .A(_04502_ ), .B1(_04544_ ), .B2(_04545_ ), .ZN(_04546_ ) );
AND2_X1 _11859_ ( .A1(_03080_ ), .A2(\u_exu.alu_p1[17] ), .ZN(_04547_ ) );
AND2_X1 _11860_ ( .A1(\u_exu.alu_p1[16] ), .A2(fanout_net_14 ), .ZN(_04548_ ) );
OAI21_X1 _11861_ ( .A(fanout_net_15 ), .B1(_04547_ ), .B2(_04548_ ), .ZN(_04549_ ) );
NAND2_X1 _11862_ ( .A1(_04546_ ), .A2(_04549_ ), .ZN(_04550_ ) );
NAND2_X1 _11863_ ( .A1(_04550_ ), .A2(fanout_net_17 ), .ZN(_04551_ ) );
AND2_X1 _11864_ ( .A1(_03080_ ), .A2(\u_exu.alu_p1[21] ), .ZN(_04552_ ) );
AND2_X1 _11865_ ( .A1(\u_exu.alu_p1[20] ), .A2(fanout_net_14 ), .ZN(_04553_ ) );
OR3_X1 _11866_ ( .A1(_04552_ ), .A2(_04483_ ), .A3(_04553_ ), .ZN(_04554_ ) );
NOR2_X1 _11867_ ( .A1(_03265_ ), .A2(fanout_net_14 ), .ZN(_04555_ ) );
INV_X1 _11868_ ( .A(_04555_ ), .ZN(_04556_ ) );
AND2_X1 _11869_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[22] ), .ZN(_04557_ ) );
INV_X1 _11870_ ( .A(_04557_ ), .ZN(_04558_ ) );
NAND3_X1 _11871_ ( .A1(_04556_ ), .A2(_04528_ ), .A3(_04558_ ), .ZN(_04559_ ) );
NAND3_X1 _11872_ ( .A1(_04554_ ), .A2(_04498_ ), .A3(_04559_ ), .ZN(_04560_ ) );
NAND3_X1 _11873_ ( .A1(_04551_ ), .A2(_04560_ ), .A3(fanout_net_19 ), .ZN(_04561_ ) );
AND2_X2 _11874_ ( .A1(_03378_ ), .A2(_03418_ ), .ZN(_04562_ ) );
CLKBUF_X2 _11875_ ( .A(_04562_ ), .Z(_04563_ ) );
NAND3_X1 _11876_ ( .A1(_04543_ ), .A2(_04561_ ), .A3(_04563_ ), .ZN(_04564_ ) );
BUF_X4 _11877_ ( .A(_03374_ ), .Z(_04565_ ) );
OAI211_X1 _11878_ ( .A(_04565_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_ctrl[0] ), .C2(\u_exu.alu_p2[31] ), .ZN(_04566_ ) );
NAND2_X1 _11879_ ( .A1(\u_exu.alu_ctrl[0] ), .A2(\u_exu.alu_p2[31] ), .ZN(_04567_ ) );
AOI21_X1 _11880_ ( .A(_04566_ ), .B1(_03361_ ), .B2(_04567_ ), .ZN(_04568_ ) );
NAND4_X1 _11881_ ( .A1(_04531_ ), .A2(_03454_ ), .A3(_03457_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B_$_MUX__B_A_$_NAND__Y_B ), .ZN(_04569_ ) );
MUX2_X1 _11882_ ( .A(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ), .B(_04569_ ), .S(_03366_ ), .Z(_04570_ ) );
BUF_X4 _11883_ ( .A(_03381_ ), .Z(_04571_ ) );
NOR2_X1 _11884_ ( .A1(_04570_ ), .A2(_04571_ ), .ZN(_04572_ ) );
BUF_X4 _11885_ ( .A(_03084_ ), .Z(_04573_ ) );
BUF_X4 _11886_ ( .A(_04573_ ), .Z(_04574_ ) );
AOI211_X1 _11887_ ( .A(_04568_ ), .B(_04572_ ), .C1(_03098_ ), .C2(_04574_ ), .ZN(_04575_ ) );
NAND4_X1 _11888_ ( .A1(_04480_ ), .A2(_04522_ ), .A3(_04564_ ), .A4(_04575_ ), .ZN(_04576_ ) );
BUF_X4 _11889_ ( .A(_03071_ ), .Z(_04577_ ) );
BUF_X4 _11890_ ( .A(_04577_ ), .Z(_04578_ ) );
MUX2_X1 _11891_ ( .A(\u_exu.alu_p1[31] ), .B(_04576_ ), .S(_04578_ ), .Z(_04579_ ) );
CLKBUF_X2 _11892_ ( .A(_01060_ ), .Z(_04580_ ) );
NAND2_X1 _11893_ ( .A1(_04579_ ), .A2(_04580_ ), .ZN(_04581_ ) );
INV_X1 _11894_ ( .A(_04581_ ), .ZN(_00303_ ) );
AOI211_X1 _11895_ ( .A(_00898_ ), .B(_04476_ ), .C1(_00745_ ), .C2(_00759_ ), .ZN(_00304_ ) );
BUF_X4 _11896_ ( .A(_00897_ ), .Z(_04582_ ) );
CLKBUF_X2 _11897_ ( .A(_03373_ ), .Z(_04583_ ) );
CLKBUF_X2 _11898_ ( .A(_03077_ ), .Z(_04584_ ) );
AND4_X1 _11899_ ( .A1(_03144_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(fanout_net_20 ), .ZN(_04585_ ) );
BUF_X4 _11900_ ( .A(_04478_ ), .Z(_04586_ ) );
NAND3_X1 _11901_ ( .A1(_03353_ ), .A2(_03146_ ), .A3(_03356_ ), .ZN(_04587_ ) );
NAND3_X1 _11902_ ( .A1(_03358_ ), .A2(_04586_ ), .A3(_04587_ ), .ZN(_04588_ ) );
AND2_X1 _11903_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[3] ), .ZN(_04589_ ) );
OR3_X1 _11904_ ( .A1(_03428_ ), .A2(_04589_ ), .A3(_04482_ ), .ZN(_04590_ ) );
OR3_X1 _11905_ ( .A1(_03425_ ), .A2(_03429_ ), .A3(fanout_net_15 ), .ZN(_04591_ ) );
AOI21_X1 _11906_ ( .A(fanout_net_17 ), .B1(_04590_ ), .B2(_04591_ ), .ZN(_04592_ ) );
NOR2_X1 _11907_ ( .A1(_03225_ ), .A2(fanout_net_14 ), .ZN(_04593_ ) );
AND2_X1 _11908_ ( .A1(fanout_net_14 ), .A2(\u_exu.alu_p1[1] ), .ZN(_04594_ ) );
OR3_X1 _11909_ ( .A1(_04593_ ), .A2(_04594_ ), .A3(fanout_net_15 ), .ZN(_04595_ ) );
OAI21_X1 _11910_ ( .A(_04595_ ), .B1(_04502_ ), .B2(_03420_ ), .ZN(_04596_ ) );
AOI21_X1 _11911_ ( .A(_04592_ ), .B1(fanout_net_17 ), .B2(_04596_ ), .ZN(_04597_ ) );
OR2_X1 _11912_ ( .A1(_04597_ ), .A2(_04523_ ), .ZN(_04598_ ) );
BUF_X2 _11913_ ( .A(_03453_ ), .Z(_04599_ ) );
BUF_X2 _11914_ ( .A(_04599_ ), .Z(_04600_ ) );
OR3_X1 _11915_ ( .A1(_03445_ ), .A2(_03426_ ), .A3(_04496_ ), .ZN(_04601_ ) );
OR3_X1 _11916_ ( .A1(_03442_ ), .A2(_03446_ ), .A3(fanout_net_15 ), .ZN(_04602_ ) );
AOI21_X1 _11917_ ( .A(_04490_ ), .B1(_04601_ ), .B2(_04602_ ), .ZN(_04603_ ) );
OR3_X1 _11918_ ( .A1(_03434_ ), .A2(_03443_ ), .A3(_04496_ ), .ZN(_04604_ ) );
OR3_X1 _11919_ ( .A1(_03437_ ), .A2(_03435_ ), .A3(fanout_net_15 ), .ZN(_04605_ ) );
AOI21_X1 _11920_ ( .A(fanout_net_17 ), .B1(_04604_ ), .B2(_04605_ ), .ZN(_04606_ ) );
OAI21_X1 _11921_ ( .A(_04600_ ), .B1(_04603_ ), .B2(_04606_ ), .ZN(_04607_ ) );
AND3_X1 _11922_ ( .A1(_04598_ ), .A2(_04501_ ), .A3(_04607_ ), .ZN(_04608_ ) );
NOR2_X1 _11923_ ( .A1(_03366_ ), .A2(\u_exu.alu_p2[4] ), .ZN(_04609_ ) );
NAND3_X1 _11924_ ( .A1(_03412_ ), .A2(_03456_ ), .A3(_04483_ ), .ZN(_04610_ ) );
OAI21_X1 _11925_ ( .A(\u_exu.alu_p1[31] ), .B1(fanout_net_17 ), .B2(fanout_net_15 ), .ZN(_04611_ ) );
AOI21_X1 _11926_ ( .A(fanout_net_19 ), .B1(_04610_ ), .B2(_04611_ ), .ZN(_04612_ ) );
AND2_X1 _11927_ ( .A1(\u_exu.alu_p1[31] ), .A2(fanout_net_19 ), .ZN(_04613_ ) );
OAI21_X1 _11928_ ( .A(_04609_ ), .B1(_04612_ ), .B2(_04613_ ), .ZN(_04614_ ) );
AND2_X2 _11929_ ( .A1(\u_exu.alu_ctrl[1] ), .A2(\u_exu.alu_p2[4] ), .ZN(_04615_ ) );
AND2_X1 _11930_ ( .A1(_04615_ ), .A2(\u_exu.alu_p1[31] ), .ZN(_04616_ ) );
NOR2_X1 _11931_ ( .A1(_04610_ ), .A2(fanout_net_19 ), .ZN(_04617_ ) );
NOR2_X1 _11932_ ( .A1(\u_exu.alu_ctrl[1] ), .A2(\u_exu.alu_p2[4] ), .ZN(_04618_ ) );
AOI21_X1 _11933_ ( .A(_04616_ ), .B1(_04617_ ), .B2(_04618_ ), .ZN(_04619_ ) );
AOI21_X1 _11934_ ( .A(_04571_ ), .B1(_04614_ ), .B2(_04619_ ), .ZN(_04620_ ) );
OR3_X1 _11935_ ( .A1(_03408_ ), .A2(_03400_ ), .A3(_04528_ ), .ZN(_04621_ ) );
MUX2_X1 _11936_ ( .A(\u_exu.alu_p1[30] ), .B(\u_exu.alu_p1[29] ), .S(fanout_net_14 ), .Z(_04622_ ) );
OAI211_X1 _11937_ ( .A(_04621_ ), .B(_04490_ ), .C1(fanout_net_15 ), .C2(_04622_ ), .ZN(_04623_ ) );
OAI211_X1 _11938_ ( .A(_03405_ ), .B(_04502_ ), .C1(\u_exu.alu_p2[0] ), .C2(_03321_ ), .ZN(_04624_ ) );
NAND3_X1 _11939_ ( .A1(_03403_ ), .A2(fanout_net_15 ), .A3(_03395_ ), .ZN(_04625_ ) );
NAND3_X1 _11940_ ( .A1(_04624_ ), .A2(_04625_ ), .A3(fanout_net_17 ), .ZN(_04626_ ) );
NAND3_X1 _11941_ ( .A1(_04623_ ), .A2(_04520_ ), .A3(_04626_ ), .ZN(_04627_ ) );
OAI21_X1 _11942_ ( .A(_04483_ ), .B1(_03382_ ), .B2(_03387_ ), .ZN(_04628_ ) );
OAI21_X1 _11943_ ( .A(fanout_net_15 ), .B1(_03386_ ), .B2(_03438_ ), .ZN(_04629_ ) );
NAND2_X1 _11944_ ( .A1(_04628_ ), .A2(_04629_ ), .ZN(_04630_ ) );
NAND2_X1 _11945_ ( .A1(_04630_ ), .A2(fanout_net_17 ), .ZN(_04631_ ) );
OR3_X1 _11946_ ( .A1(_03391_ ), .A2(_03383_ ), .A3(_04483_ ), .ZN(_04632_ ) );
NOR2_X1 _11947_ ( .A1(_03269_ ), .A2(\u_exu.alu_p2[0] ), .ZN(_04633_ ) );
OR3_X1 _11948_ ( .A1(_04633_ ), .A2(_03392_ ), .A3(fanout_net_15 ), .ZN(_04634_ ) );
NAND3_X1 _11949_ ( .A1(_04632_ ), .A2(_04634_ ), .A3(_04490_ ), .ZN(_04635_ ) );
NAND3_X1 _11950_ ( .A1(_04631_ ), .A2(_04635_ ), .A3(fanout_net_19 ), .ZN(_04636_ ) );
BUF_X2 _11951_ ( .A(_04562_ ), .Z(_04637_ ) );
AND3_X1 _11952_ ( .A1(_04627_ ), .A2(_04636_ ), .A3(_04637_ ), .ZN(_04638_ ) );
BUF_X2 _11953_ ( .A(_04573_ ), .Z(_04639_ ) );
NAND2_X1 _11954_ ( .A1(_03125_ ), .A2(_04639_ ), .ZN(_04640_ ) );
AOI21_X1 _11955_ ( .A(\u_exu.alu_p1[30] ), .B1(\u_exu.alu_ctrl[0] ), .B2(\u_exu.alu_p2[30] ), .ZN(_04641_ ) );
BUF_X4 _11956_ ( .A(_04565_ ), .Z(_04642_ ) );
OAI211_X1 _11957_ ( .A(_04642_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_ctrl[0] ), .C2(\u_exu.alu_p2[30] ), .ZN(_04643_ ) );
OAI211_X1 _11958_ ( .A(_04640_ ), .B(_03071_ ), .C1(_04641_ ), .C2(_04643_ ), .ZN(_04644_ ) );
NOR4_X1 _11959_ ( .A1(_04608_ ), .A2(_04620_ ), .A3(_04638_ ), .A4(_04644_ ), .ZN(_04645_ ) );
AOI211_X1 _11960_ ( .A(_04582_ ), .B(_04585_ ), .C1(_04588_ ), .C2(_04645_ ), .ZN(_00305_ ) );
NOR4_X1 _11961_ ( .A1(_03379_ ), .A2(\u_exu.alu_p1[21] ), .A3(\u_exu.alu_ctrl[5] ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_04646_ ) );
NAND2_X1 _11962_ ( .A1(_03254_ ), .A2(_03287_ ), .ZN(_04647_ ) );
AND2_X1 _11963_ ( .A1(_04647_ ), .A2(_03299_ ), .ZN(_04648_ ) );
NOR2_X1 _11964_ ( .A1(_03256_ ), .A2(\u_exu.alu_p1[20] ), .ZN(_04649_ ) );
NOR3_X1 _11965_ ( .A1(_04648_ ), .A2(_03304_ ), .A3(_04649_ ), .ZN(_04650_ ) );
OR3_X1 _11966_ ( .A1(_04650_ ), .A2(_03261_ ), .A3(_03304_ ), .ZN(_04651_ ) );
OAI21_X1 _11967_ ( .A(_03261_ ), .B1(_04650_ ), .B2(_03304_ ), .ZN(_04652_ ) );
NAND3_X1 _11968_ ( .A1(_04651_ ), .A2(_04586_ ), .A3(_04652_ ), .ZN(_04653_ ) );
NOR2_X1 _11969_ ( .A1(_04537_ ), .A2(_04534_ ), .ZN(_04654_ ) );
NOR2_X1 _11970_ ( .A1(_03317_ ), .A2(\u_exu.alu_p2[0] ), .ZN(_04655_ ) );
NOR2_X1 _11971_ ( .A1(_04655_ ), .A2(_04526_ ), .ZN(_04656_ ) );
MUX2_X1 _11972_ ( .A(_04654_ ), .B(_04656_ ), .S(fanout_net_15 ), .Z(_04657_ ) );
NAND2_X1 _11973_ ( .A1(_04657_ ), .A2(fanout_net_17 ), .ZN(_04658_ ) );
CLKBUF_X2 _11974_ ( .A(_03413_ ), .Z(_04659_ ) );
OAI21_X1 _11975_ ( .A(_04659_ ), .B1(_04552_ ), .B2(_04557_ ), .ZN(_04660_ ) );
OAI21_X1 _11976_ ( .A(fanout_net_15 ), .B1(_04555_ ), .B2(_04539_ ), .ZN(_04661_ ) );
NAND2_X1 _11977_ ( .A1(_04660_ ), .A2(_04661_ ), .ZN(_04662_ ) );
OAI21_X1 _11978_ ( .A(_04658_ ), .B1(fanout_net_17 ), .B2(_04662_ ), .ZN(_04663_ ) );
NOR2_X1 _11979_ ( .A1(_04663_ ), .A2(fanout_net_19 ), .ZN(_04664_ ) );
AND2_X1 _11980_ ( .A1(\u_exu.alu_p1[31] ), .A2(fanout_net_17 ), .ZN(_04665_ ) );
MUX2_X1 _11981_ ( .A(_03347_ ), .B(_03144_ ), .S(\u_exu.alu_p2[0] ), .Z(_04666_ ) );
INV_X1 _11982_ ( .A(_04666_ ), .ZN(_04667_ ) );
MUX2_X1 _11983_ ( .A(\u_exu.alu_p1[31] ), .B(_04667_ ), .S(_04482_ ), .Z(_04668_ ) );
AOI21_X1 _11984_ ( .A(_04665_ ), .B1(_04668_ ), .B2(_03456_ ), .ZN(_04669_ ) );
NOR2_X1 _11985_ ( .A1(_04669_ ), .A2(_04518_ ), .ZN(_04670_ ) );
OAI21_X1 _11986_ ( .A(_04609_ ), .B1(_04664_ ), .B2(_04670_ ), .ZN(_04671_ ) );
AND3_X1 _11987_ ( .A1(_03080_ ), .A2(\u_exu.alu_p1[31] ), .A3(fanout_net_15 ), .ZN(_04672_ ) );
AOI21_X1 _11988_ ( .A(_04672_ ), .B1(_04667_ ), .B2(_04496_ ), .ZN(_04673_ ) );
NOR3_X1 _11989_ ( .A1(_04673_ ), .A2(_03453_ ), .A3(fanout_net_17 ), .ZN(_04674_ ) );
OAI21_X1 _11990_ ( .A(_04618_ ), .B1(_04664_ ), .B2(_04674_ ), .ZN(_04675_ ) );
AND2_X1 _11991_ ( .A1(_04671_ ), .A2(_04675_ ), .ZN(_04676_ ) );
INV_X1 _11992_ ( .A(_04616_ ), .ZN(_04677_ ) );
AOI21_X1 _11993_ ( .A(_04571_ ), .B1(_04676_ ), .B2(_04677_ ), .ZN(_04678_ ) );
BUF_X4 _11994_ ( .A(_03418_ ), .Z(_04679_ ) );
OAI21_X1 _11995_ ( .A(_04502_ ), .B1(_04506_ ), .B2(_04507_ ), .ZN(_04680_ ) );
OAI21_X1 _11996_ ( .A(fanout_net_15 ), .B1(_04486_ ), .B2(_04487_ ), .ZN(_04681_ ) );
NAND2_X1 _11997_ ( .A1(_04680_ ), .A2(_04681_ ), .ZN(_04682_ ) );
NAND2_X1 _11998_ ( .A1(_04682_ ), .A2(fanout_net_17 ), .ZN(_04683_ ) );
OAI21_X1 _11999_ ( .A(fanout_net_15 ), .B1(_04503_ ), .B2(_04504_ ), .ZN(_04684_ ) );
OAI21_X1 _12000_ ( .A(_04502_ ), .B1(_04514_ ), .B2(_04515_ ), .ZN(_04685_ ) );
NAND2_X1 _12001_ ( .A1(_04684_ ), .A2(_04685_ ), .ZN(_04686_ ) );
NAND2_X1 _12002_ ( .A1(_04686_ ), .A2(_04490_ ), .ZN(_04687_ ) );
NAND2_X1 _12003_ ( .A1(_04683_ ), .A2(_04687_ ), .ZN(_04688_ ) );
OAI21_X1 _12004_ ( .A(_04679_ ), .B1(_04688_ ), .B2(_04524_ ), .ZN(_04689_ ) );
INV_X1 _12005_ ( .A(_03378_ ), .ZN(_04690_ ) );
OAI21_X1 _12006_ ( .A(_04502_ ), .B1(_04547_ ), .B2(_04548_ ), .ZN(_04691_ ) );
OAI21_X1 _12007_ ( .A(fanout_net_16 ), .B1(_04511_ ), .B2(_04512_ ), .ZN(_04692_ ) );
NAND2_X1 _12008_ ( .A1(_04691_ ), .A2(_04692_ ), .ZN(_04693_ ) );
NAND2_X1 _12009_ ( .A1(_04693_ ), .A2(fanout_net_17 ), .ZN(_04694_ ) );
OR3_X1 _12010_ ( .A1(_04544_ ), .A2(_04483_ ), .A3(_04545_ ), .ZN(_04695_ ) );
OR3_X1 _12011_ ( .A1(_04552_ ), .A2(fanout_net_16 ), .A3(_04553_ ), .ZN(_04696_ ) );
NAND3_X1 _12012_ ( .A1(_04695_ ), .A2(_04696_ ), .A3(_04490_ ), .ZN(_04697_ ) );
AND3_X1 _12013_ ( .A1(_04694_ ), .A2(_04697_ ), .A3(_04600_ ), .ZN(_04698_ ) );
NOR3_X1 _12014_ ( .A1(_04689_ ), .A2(_04690_ ), .A3(_04698_ ), .ZN(_04699_ ) );
NAND2_X1 _12015_ ( .A1(_03080_ ), .A2(\u_exu.alu_p1[1] ), .ZN(_04700_ ) );
AOI21_X1 _12016_ ( .A(fanout_net_16 ), .B1(_03464_ ), .B2(_04700_ ), .ZN(_04701_ ) );
OAI21_X1 _12017_ ( .A(_04496_ ), .B1(_04481_ ), .B2(_04484_ ), .ZN(_04702_ ) );
OAI21_X1 _12018_ ( .A(fanout_net_16 ), .B1(_04493_ ), .B2(_04494_ ), .ZN(_04703_ ) );
NAND2_X1 _12019_ ( .A1(_04702_ ), .A2(_04703_ ), .ZN(_04704_ ) );
MUX2_X1 _12020_ ( .A(_04701_ ), .B(_04704_ ), .S(_03456_ ), .Z(_04705_ ) );
NAND3_X1 _12021_ ( .A1(_04705_ ), .A2(_04520_ ), .A3(_04501_ ), .ZN(_04706_ ) );
NAND2_X1 _12022_ ( .A1(_03122_ ), .A2(_04639_ ), .ZN(_04707_ ) );
AOI21_X1 _12023_ ( .A(\u_exu.alu_p1[21] ), .B1(\u_exu.alu_p2[21] ), .B2(\u_exu.alu_ctrl[0] ), .ZN(_04708_ ) );
OAI211_X1 _12024_ ( .A(_04642_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p2[21] ), .C2(\u_exu.alu_ctrl[0] ), .ZN(_04709_ ) );
OAI211_X1 _12025_ ( .A(_04706_ ), .B(_04707_ ), .C1(_04708_ ), .C2(_04709_ ), .ZN(_04710_ ) );
NOR4_X1 _12026_ ( .A1(_04678_ ), .A2(_03070_ ), .A3(_04699_ ), .A4(_04710_ ), .ZN(_04711_ ) );
AOI211_X1 _12027_ ( .A(_04582_ ), .B(_04646_ ), .C1(_04653_ ), .C2(_04711_ ), .ZN(_00306_ ) );
INV_X1 _12028_ ( .A(_04477_ ), .ZN(_04712_ ) );
CLKBUF_X2 _12029_ ( .A(_04712_ ), .Z(_04713_ ) );
INV_X1 _12030_ ( .A(_04648_ ), .ZN(_04714_ ) );
AOI21_X1 _12031_ ( .A(_04713_ ), .B1(_04714_ ), .B2(_03258_ ), .ZN(_04715_ ) );
OAI21_X1 _12032_ ( .A(_04715_ ), .B1(_03258_ ), .B2(_04714_ ), .ZN(_04716_ ) );
BUF_X4 _12033_ ( .A(_03380_ ), .Z(_04717_ ) );
INV_X1 _12034_ ( .A(_04665_ ), .ZN(_04718_ ) );
OAI21_X1 _12035_ ( .A(_04718_ ), .B1(_03414_ ), .B2(fanout_net_17 ), .ZN(_04719_ ) );
AND2_X1 _12036_ ( .A1(_04719_ ), .A2(fanout_net_19 ), .ZN(_04720_ ) );
AOI21_X1 _12037_ ( .A(fanout_net_17 ), .B1(_03393_ ), .B2(_03396_ ), .ZN(_04721_ ) );
AOI21_X1 _12038_ ( .A(_03455_ ), .B1(_03401_ ), .B2(_03406_ ), .ZN(_04722_ ) );
NOR3_X1 _12039_ ( .A1(_04721_ ), .A2(_04722_ ), .A3(fanout_net_19 ), .ZN(_04723_ ) );
OAI21_X1 _12040_ ( .A(_04609_ ), .B1(_04720_ ), .B2(_04723_ ), .ZN(_04724_ ) );
NOR3_X1 _12041_ ( .A1(_03414_ ), .A2(_04518_ ), .A3(fanout_net_17 ), .ZN(_04725_ ) );
OAI21_X1 _12042_ ( .A(_04618_ ), .B1(_04723_ ), .B2(_04725_ ), .ZN(_04726_ ) );
NAND2_X1 _12043_ ( .A1(_04724_ ), .A2(_04726_ ), .ZN(_04727_ ) );
OAI21_X1 _12044_ ( .A(_04717_ ), .B1(_04727_ ), .B2(_04616_ ), .ZN(_04728_ ) );
OAI21_X1 _12045_ ( .A(_04659_ ), .B1(_03434_ ), .B2(_03443_ ), .ZN(_04729_ ) );
OAI21_X1 _12046_ ( .A(fanout_net_16 ), .B1(_03442_ ), .B2(_03446_ ), .ZN(_04730_ ) );
AOI21_X1 _12047_ ( .A(fanout_net_17 ), .B1(_04729_ ), .B2(_04730_ ), .ZN(_04731_ ) );
OAI21_X1 _12048_ ( .A(_04659_ ), .B1(_03445_ ), .B2(_03426_ ), .ZN(_04732_ ) );
OAI21_X1 _12049_ ( .A(fanout_net_16 ), .B1(_03425_ ), .B2(_03429_ ), .ZN(_04733_ ) );
AOI21_X1 _12050_ ( .A(_03455_ ), .B1(_04732_ ), .B2(_04733_ ), .ZN(_04734_ ) );
NOR2_X1 _12051_ ( .A1(_04731_ ), .A2(_04734_ ), .ZN(_04735_ ) );
NAND2_X1 _12052_ ( .A1(_04735_ ), .A2(fanout_net_19 ), .ZN(_04736_ ) );
OAI21_X1 _12053_ ( .A(_04483_ ), .B1(_03391_ ), .B2(_03383_ ), .ZN(_04737_ ) );
OAI21_X1 _12054_ ( .A(fanout_net_16 ), .B1(_03382_ ), .B2(_03387_ ), .ZN(_04738_ ) );
NAND2_X1 _12055_ ( .A1(_04737_ ), .A2(_04738_ ), .ZN(_04739_ ) );
NAND2_X1 _12056_ ( .A1(_04739_ ), .A2(_04490_ ), .ZN(_04740_ ) );
OR3_X1 _12057_ ( .A1(_03437_ ), .A2(_03435_ ), .A3(_04496_ ), .ZN(_04741_ ) );
OR3_X1 _12058_ ( .A1(_03386_ ), .A2(_03438_ ), .A3(fanout_net_16 ), .ZN(_04742_ ) );
NAND3_X1 _12059_ ( .A1(_04741_ ), .A2(_04742_ ), .A3(fanout_net_17 ), .ZN(_04743_ ) );
NAND3_X1 _12060_ ( .A1(_04740_ ), .A2(_04743_ ), .A3(_04524_ ), .ZN(_04744_ ) );
NAND3_X1 _12061_ ( .A1(_04736_ ), .A2(_04563_ ), .A3(_04744_ ), .ZN(_04745_ ) );
OAI211_X1 _12062_ ( .A(_04642_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[20] ), .C2(\u_exu.alu_p2[20] ), .ZN(_04746_ ) );
AOI21_X1 _12063_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[20] ), .B2(\u_exu.alu_p2[20] ), .ZN(_04747_ ) );
NOR2_X1 _12064_ ( .A1(_04746_ ), .A2(_04747_ ), .ZN(_04748_ ) );
OAI21_X1 _12065_ ( .A(_03413_ ), .B1(_03428_ ), .B2(_04589_ ), .ZN(_04749_ ) );
OAI21_X1 _12066_ ( .A(fanout_net_16 ), .B1(_04593_ ), .B2(_04594_ ), .ZN(_04750_ ) );
NAND2_X1 _12067_ ( .A1(_04749_ ), .A2(_04750_ ), .ZN(_04751_ ) );
MUX2_X1 _12068_ ( .A(_03421_ ), .B(_04751_ ), .S(_03455_ ), .Z(_04752_ ) );
AND3_X1 _12069_ ( .A1(_04752_ ), .A2(_04600_ ), .A3(_04500_ ), .ZN(_04753_ ) );
AOI211_X1 _12070_ ( .A(_04748_ ), .B(_04753_ ), .C1(_03102_ ), .C2(_04574_ ), .ZN(_04754_ ) );
NAND4_X1 _12071_ ( .A1(_04716_ ), .A2(_04728_ ), .A3(_04745_ ), .A4(_04754_ ), .ZN(_04755_ ) );
MUX2_X1 _12072_ ( .A(\u_exu.alu_p1[20] ), .B(_04755_ ), .S(_04578_ ), .Z(_04756_ ) );
AND2_X1 _12073_ ( .A1(_04756_ ), .A2(_04580_ ), .ZN(_00307_ ) );
NOR4_X1 _12074_ ( .A1(_03379_ ), .A2(\u_exu.alu_p1[19] ), .A3(\u_exu.alu_ctrl[5] ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_04757_ ) );
INV_X1 _12075_ ( .A(_03275_ ), .ZN(_04758_ ) );
INV_X1 _12076_ ( .A(_03283_ ), .ZN(_04759_ ) );
AOI21_X1 _12077_ ( .A(_04759_ ), .B1(_03200_ ), .B2(_03252_ ), .ZN(_04760_ ) );
NAND2_X1 _12078_ ( .A1(_04760_ ), .A2(_03286_ ), .ZN(_04761_ ) );
AOI21_X1 _12079_ ( .A(_04758_ ), .B1(_04761_ ), .B2(_03296_ ), .ZN(_04762_ ) );
OR3_X1 _12080_ ( .A1(_04762_ ), .A2(_03278_ ), .A3(_03289_ ), .ZN(_04763_ ) );
OAI21_X1 _12081_ ( .A(_03278_ ), .B1(_04762_ ), .B2(_03289_ ), .ZN(_04764_ ) );
NAND3_X1 _12082_ ( .A1(_04763_ ), .A2(_04586_ ), .A3(_04764_ ), .ZN(_04765_ ) );
MUX2_X1 _12083_ ( .A(_04656_ ), .B(_04666_ ), .S(fanout_net_16 ), .Z(_04766_ ) );
OR2_X1 _12084_ ( .A1(_04766_ ), .A2(fanout_net_18 ), .ZN(_04767_ ) );
AOI21_X1 _12085_ ( .A(_04518_ ), .B1(_04767_ ), .B2(_04718_ ), .ZN(_04768_ ) );
OR3_X1 _12086_ ( .A1(_04552_ ), .A2(_04482_ ), .A3(_04557_ ), .ZN(_04769_ ) );
OR3_X1 _12087_ ( .A1(_04544_ ), .A2(fanout_net_16 ), .A3(_04553_ ), .ZN(_04770_ ) );
NAND3_X1 _12088_ ( .A1(_04769_ ), .A2(_04770_ ), .A3(_03455_ ), .ZN(_04771_ ) );
NAND3_X1 _12089_ ( .A1(_04538_ ), .A2(fanout_net_16 ), .A3(_04535_ ), .ZN(_04772_ ) );
NAND3_X1 _12090_ ( .A1(_04556_ ), .A2(_04496_ ), .A3(_04540_ ), .ZN(_04773_ ) );
NAND3_X1 _12091_ ( .A1(_04772_ ), .A2(_04773_ ), .A3(fanout_net_18 ), .ZN(_04774_ ) );
AOI21_X1 _12092_ ( .A(fanout_net_19 ), .B1(_04771_ ), .B2(_04774_ ), .ZN(_04775_ ) );
OAI21_X1 _12093_ ( .A(_04609_ ), .B1(_04768_ ), .B2(_04775_ ), .ZN(_04776_ ) );
NAND4_X1 _12094_ ( .A1(_04496_ ), .A2(_03080_ ), .A3(\u_exu.alu_p1[31] ), .A4(fanout_net_18 ), .ZN(_04777_ ) );
OAI21_X1 _12095_ ( .A(_04777_ ), .B1(_04766_ ), .B2(fanout_net_18 ), .ZN(_04778_ ) );
AND2_X1 _12096_ ( .A1(_04778_ ), .A2(fanout_net_19 ), .ZN(_04779_ ) );
OAI21_X1 _12097_ ( .A(_04618_ ), .B1(_04779_ ), .B2(_04775_ ), .ZN(_04780_ ) );
NAND2_X1 _12098_ ( .A1(_04776_ ), .A2(_04780_ ), .ZN(_04781_ ) );
OAI21_X1 _12099_ ( .A(_04717_ ), .B1(_04781_ ), .B2(_04616_ ), .ZN(_04782_ ) );
NAND2_X1 _12100_ ( .A1(_04509_ ), .A2(_03457_ ), .ZN(_04783_ ) );
NAND3_X1 _12101_ ( .A1(_04485_ ), .A2(_04488_ ), .A3(fanout_net_18 ), .ZN(_04784_ ) );
NAND3_X1 _12102_ ( .A1(_04783_ ), .A2(_04784_ ), .A3(fanout_net_19 ), .ZN(_04785_ ) );
NAND2_X1 _12103_ ( .A1(_04550_ ), .A2(_03457_ ), .ZN(_04786_ ) );
NAND3_X1 _12104_ ( .A1(_04513_ ), .A2(fanout_net_18 ), .A3(_04516_ ), .ZN(_04787_ ) );
NAND3_X1 _12105_ ( .A1(_04786_ ), .A2(_04787_ ), .A3(_04600_ ), .ZN(_04788_ ) );
NAND3_X1 _12106_ ( .A1(_04785_ ), .A2(_04788_ ), .A3(_04637_ ), .ZN(_04789_ ) );
NOR2_X1 _12107_ ( .A1(_04497_ ), .A2(fanout_net_18 ), .ZN(_04790_ ) );
NAND3_X1 _12108_ ( .A1(_04790_ ), .A2(_04524_ ), .A3(_04501_ ), .ZN(_04791_ ) );
OAI211_X1 _12109_ ( .A(_04565_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[19] ), .C2(\u_exu.alu_p2[19] ), .ZN(_04792_ ) );
AOI21_X1 _12110_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[19] ), .B2(\u_exu.alu_p2[19] ), .ZN(_04793_ ) );
NOR2_X1 _12111_ ( .A1(_04792_ ), .A2(_04793_ ), .ZN(_04794_ ) );
AOI211_X1 _12112_ ( .A(_03070_ ), .B(_04794_ ), .C1(_03103_ ), .C2(_04639_ ), .ZN(_04795_ ) );
AND4_X1 _12113_ ( .A1(_04782_ ), .A2(_04789_ ), .A3(_04791_ ), .A4(_04795_ ), .ZN(_04796_ ) );
AOI211_X1 _12114_ ( .A(_04582_ ), .B(_04757_ ), .C1(_04765_ ), .C2(_04796_ ), .ZN(_00308_ ) );
AND4_X1 _12115_ ( .A1(_03274_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(fanout_net_20 ), .ZN(_04797_ ) );
AOI211_X1 _12116_ ( .A(_03275_ ), .B(_03297_ ), .C1(_04760_ ), .C2(_03286_ ), .ZN(_04798_ ) );
OR3_X1 _12117_ ( .A1(_04762_ ), .A2(_04798_ ), .A3(_04713_ ), .ZN(_04799_ ) );
AOI21_X1 _12118_ ( .A(_04489_ ), .B1(_04590_ ), .B2(_04591_ ), .ZN(_04800_ ) );
AOI21_X1 _12119_ ( .A(fanout_net_18 ), .B1(_04601_ ), .B2(_04602_ ), .ZN(_04801_ ) );
OAI21_X1 _12120_ ( .A(fanout_net_19 ), .B1(_04800_ ), .B2(_04801_ ), .ZN(_04802_ ) );
AOI21_X1 _12121_ ( .A(_04489_ ), .B1(_04604_ ), .B2(_04605_ ), .ZN(_04803_ ) );
AND3_X1 _12122_ ( .A1(_04628_ ), .A2(_04629_ ), .A3(_03456_ ), .ZN(_04804_ ) );
OAI21_X1 _12123_ ( .A(_04523_ ), .B1(_04803_ ), .B2(_04804_ ), .ZN(_04805_ ) );
AND3_X1 _12124_ ( .A1(_04802_ ), .A2(_04637_ ), .A3(_04805_ ), .ZN(_04806_ ) );
NOR2_X1 _12125_ ( .A1(_04596_ ), .A2(fanout_net_18 ), .ZN(_04807_ ) );
NAND3_X1 _12126_ ( .A1(_04807_ ), .A2(_04600_ ), .A3(_04501_ ), .ZN(_04808_ ) );
OAI211_X1 _12127_ ( .A(_03374_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[18] ), .C2(\u_exu.alu_p2[18] ), .ZN(_04809_ ) );
AOI21_X1 _12128_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[18] ), .B2(\u_exu.alu_p2[18] ), .ZN(_04810_ ) );
OR2_X1 _12129_ ( .A1(_04809_ ), .A2(_04810_ ), .ZN(_04811_ ) );
NAND2_X1 _12130_ ( .A1(_03121_ ), .A2(_04573_ ), .ZN(_04812_ ) );
NAND4_X1 _12131_ ( .A1(_04808_ ), .A2(_03071_ ), .A3(_04811_ ), .A4(_04812_ ), .ZN(_04813_ ) );
NAND3_X1 _12132_ ( .A1(_03412_ ), .A2(fanout_net_18 ), .A3(_04659_ ), .ZN(_04814_ ) );
OAI21_X1 _12133_ ( .A(_03413_ ), .B1(_03399_ ), .B2(_03400_ ), .ZN(_04815_ ) );
OAI21_X1 _12134_ ( .A(fanout_net_16 ), .B1(_03408_ ), .B2(_03409_ ), .ZN(_04816_ ) );
AND2_X1 _12135_ ( .A1(_04815_ ), .A2(_04816_ ), .ZN(_04817_ ) );
OAI21_X1 _12136_ ( .A(_04814_ ), .B1(_04817_ ), .B2(fanout_net_18 ), .ZN(_04818_ ) );
AND3_X1 _12137_ ( .A1(\u_exu.alu_p1[31] ), .A2(fanout_net_18 ), .A3(fanout_net_16 ), .ZN(_04819_ ) );
NOR2_X1 _12138_ ( .A1(_04818_ ), .A2(_04819_ ), .ZN(_04820_ ) );
NOR2_X1 _12139_ ( .A1(_04820_ ), .A2(_04523_ ), .ZN(_04821_ ) );
OR3_X1 _12140_ ( .A1(_03391_ ), .A2(_03392_ ), .A3(_04659_ ), .ZN(_04822_ ) );
OR3_X1 _12141_ ( .A1(_03382_ ), .A2(_03383_ ), .A3(fanout_net_16 ), .ZN(_04823_ ) );
AOI21_X1 _12142_ ( .A(fanout_net_18 ), .B1(_04822_ ), .B2(_04823_ ), .ZN(_04824_ ) );
OAI21_X1 _12143_ ( .A(_04482_ ), .B1(_04633_ ), .B2(_03394_ ), .ZN(_04825_ ) );
OAI21_X1 _12144_ ( .A(fanout_net_16 ), .B1(_03402_ ), .B2(_03404_ ), .ZN(_04826_ ) );
AND3_X1 _12145_ ( .A1(_04825_ ), .A2(_04826_ ), .A3(fanout_net_18 ), .ZN(_04827_ ) );
NOR3_X1 _12146_ ( .A1(_04824_ ), .A2(_04827_ ), .A3(fanout_net_19 ), .ZN(_04828_ ) );
OAI21_X1 _12147_ ( .A(_04609_ ), .B1(_04821_ ), .B2(_04828_ ), .ZN(_04829_ ) );
AND2_X1 _12148_ ( .A1(_04818_ ), .A2(fanout_net_19 ), .ZN(_04830_ ) );
OAI21_X1 _12149_ ( .A(_04618_ ), .B1(_04830_ ), .B2(_04828_ ), .ZN(_04831_ ) );
NAND3_X1 _12150_ ( .A1(_04829_ ), .A2(_04677_ ), .A3(_04831_ ), .ZN(_04832_ ) );
AOI211_X1 _12151_ ( .A(_04806_ ), .B(_04813_ ), .C1(_04832_ ), .C2(_04717_ ), .ZN(_04833_ ) );
AOI211_X1 _12152_ ( .A(_04582_ ), .B(_04797_ ), .C1(_04799_ ), .C2(_04833_ ), .ZN(_00309_ ) );
NOR4_X1 _12153_ ( .A1(_03379_ ), .A2(\u_exu.alu_p1[17] ), .A3(\u_exu.alu_ctrl[5] ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_04834_ ) );
OR3_X1 _12154_ ( .A1(_04760_ ), .A2(_03295_ ), .A3(_03286_ ), .ZN(_04835_ ) );
OAI21_X1 _12155_ ( .A(_03286_ ), .B1(_04760_ ), .B2(_03295_ ), .ZN(_04836_ ) );
NAND3_X1 _12156_ ( .A1(_04835_ ), .A2(_04586_ ), .A3(_04836_ ), .ZN(_04837_ ) );
MUX2_X1 _12157_ ( .A(_04673_ ), .B(_04657_ ), .S(_03456_ ), .Z(_04838_ ) );
NOR2_X1 _12158_ ( .A1(_04838_ ), .A2(_04599_ ), .ZN(_04839_ ) );
OR3_X1 _12159_ ( .A1(_04544_ ), .A2(_04659_ ), .A3(_04553_ ), .ZN(_04840_ ) );
OR3_X1 _12160_ ( .A1(_04547_ ), .A2(fanout_net_16 ), .A3(_04545_ ), .ZN(_04841_ ) );
NAND3_X1 _12161_ ( .A1(_04840_ ), .A2(_04841_ ), .A3(_04489_ ), .ZN(_04842_ ) );
NAND2_X1 _12162_ ( .A1(_04662_ ), .A2(fanout_net_18 ), .ZN(_04843_ ) );
AOI21_X1 _12163_ ( .A(fanout_net_19 ), .B1(_04842_ ), .B2(_04843_ ), .ZN(_04844_ ) );
OAI21_X1 _12164_ ( .A(_04618_ ), .B1(_04839_ ), .B2(_04844_ ), .ZN(_04845_ ) );
AND2_X1 _12165_ ( .A1(_04845_ ), .A2(_04677_ ), .ZN(_04846_ ) );
NOR2_X1 _12166_ ( .A1(_04657_ ), .A2(fanout_net_18 ), .ZN(_04847_ ) );
AOI21_X1 _12167_ ( .A(_04847_ ), .B1(fanout_net_18 ), .B2(_04668_ ), .ZN(_04848_ ) );
NOR2_X1 _12168_ ( .A1(_04848_ ), .A2(_04523_ ), .ZN(_04849_ ) );
OAI21_X1 _12169_ ( .A(_04609_ ), .B1(_04849_ ), .B2(_04844_ ), .ZN(_04850_ ) );
AOI21_X1 _12170_ ( .A(_04571_ ), .B1(_04846_ ), .B2(_04850_ ), .ZN(_04851_ ) );
NAND2_X1 _12171_ ( .A1(_04693_ ), .A2(_03457_ ), .ZN(_04852_ ) );
NAND2_X1 _12172_ ( .A1(_04686_ ), .A2(fanout_net_18 ), .ZN(_04853_ ) );
NAND3_X1 _12173_ ( .A1(_04852_ ), .A2(_04853_ ), .A3(_04519_ ), .ZN(_04854_ ) );
NAND2_X1 _12174_ ( .A1(_04854_ ), .A2(_04637_ ), .ZN(_04855_ ) );
NAND3_X1 _12175_ ( .A1(_04702_ ), .A2(_04703_ ), .A3(fanout_net_18 ), .ZN(_04856_ ) );
NAND3_X1 _12176_ ( .A1(_04680_ ), .A2(_04681_ ), .A3(_04489_ ), .ZN(_04857_ ) );
NAND2_X1 _12177_ ( .A1(_04856_ ), .A2(_04857_ ), .ZN(_04858_ ) );
AOI21_X1 _12178_ ( .A(_04855_ ), .B1(fanout_net_19 ), .B2(_04858_ ), .ZN(_04859_ ) );
NOR3_X1 _12179_ ( .A1(_04492_ ), .A2(fanout_net_18 ), .A3(fanout_net_16 ), .ZN(_04860_ ) );
AND3_X1 _12180_ ( .A1(_04860_ ), .A2(_04600_ ), .A3(_04500_ ), .ZN(_04861_ ) );
NAND2_X1 _12181_ ( .A1(_03120_ ), .A2(_04573_ ), .ZN(_04862_ ) );
AOI21_X1 _12182_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p2[17] ), .B2(\u_exu.alu_p1[17] ), .ZN(_04863_ ) );
OAI211_X1 _12183_ ( .A(_04565_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p2[17] ), .C2(\u_exu.alu_p1[17] ), .ZN(_04864_ ) );
OAI211_X1 _12184_ ( .A(_04862_ ), .B(_03071_ ), .C1(_04863_ ), .C2(_04864_ ), .ZN(_04865_ ) );
NOR4_X1 _12185_ ( .A1(_04851_ ), .A2(_04859_ ), .A3(_04861_ ), .A4(_04865_ ), .ZN(_04866_ ) );
AOI211_X1 _12186_ ( .A(_04582_ ), .B(_04834_ ), .C1(_04837_ ), .C2(_04866_ ), .ZN(_00310_ ) );
AND4_X1 _12187_ ( .A1(_03282_ ), .A2(_03373_ ), .A3(_03077_ ), .A4(fanout_net_20 ), .ZN(_04867_ ) );
OAI21_X1 _12188_ ( .A(_04478_ ), .B1(_03253_ ), .B2(_04759_ ), .ZN(_04868_ ) );
AOI21_X1 _12189_ ( .A(_04868_ ), .B1(_03253_ ), .B2(_04759_ ), .ZN(_04869_ ) );
INV_X1 _12190_ ( .A(_04637_ ), .ZN(_04870_ ) );
AOI21_X1 _12191_ ( .A(fanout_net_18 ), .B1(_04741_ ), .B2(_04742_ ), .ZN(_04871_ ) );
AND3_X1 _12192_ ( .A1(_04729_ ), .A2(_04730_ ), .A3(fanout_net_18 ), .ZN(_04872_ ) );
OR3_X1 _12193_ ( .A1(_04871_ ), .A2(_04872_ ), .A3(fanout_net_19 ), .ZN(_04873_ ) );
NAND3_X1 _12194_ ( .A1(_04749_ ), .A2(_04750_ ), .A3(fanout_net_18 ), .ZN(_04874_ ) );
NAND3_X1 _12195_ ( .A1(_04732_ ), .A2(_04733_ ), .A3(_04489_ ), .ZN(_04875_ ) );
NAND3_X1 _12196_ ( .A1(_04874_ ), .A2(_04875_ ), .A3(fanout_net_19 ), .ZN(_04876_ ) );
AOI21_X1 _12197_ ( .A(_04870_ ), .B1(_04873_ ), .B2(_04876_ ), .ZN(_04877_ ) );
AND3_X1 _12198_ ( .A1(_03420_ ), .A2(_04490_ ), .A3(_04528_ ), .ZN(_04878_ ) );
AND3_X1 _12199_ ( .A1(_04501_ ), .A2(_04600_ ), .A3(_04878_ ), .ZN(_04879_ ) );
OR4_X1 _12200_ ( .A1(_03379_ ), .A2(_03105_ ), .A3(_03373_ ), .A4(_03077_ ), .ZN(_04880_ ) );
OAI211_X1 _12201_ ( .A(_04642_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_ctrl[0] ), .C2(_03105_ ), .ZN(_04881_ ) );
AOI21_X1 _12202_ ( .A(_03106_ ), .B1(_04880_ ), .B2(_04881_ ), .ZN(_04882_ ) );
NOR4_X1 _12203_ ( .A1(_04869_ ), .A2(_04877_ ), .A3(_04879_ ), .A4(_04882_ ), .ZN(_04883_ ) );
NAND2_X1 _12204_ ( .A1(_03416_ ), .A2(_04679_ ), .ZN(_04884_ ) );
AOI21_X1 _12205_ ( .A(_04571_ ), .B1(_04884_ ), .B2(_04677_ ), .ZN(_04885_ ) );
NOR2_X1 _12206_ ( .A1(_04885_ ), .A2(_03070_ ), .ZN(_04886_ ) );
AOI211_X1 _12207_ ( .A(_04582_ ), .B(_04867_ ), .C1(_04883_ ), .C2(_04886_ ), .ZN(_00311_ ) );
NOR4_X1 _12208_ ( .A1(_03379_ ), .A2(\u_exu.alu_p1[15] ), .A3(\u_exu.alu_ctrl[5] ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_04887_ ) );
INV_X1 _12209_ ( .A(_03180_ ), .ZN(_04888_ ) );
INV_X1 _12210_ ( .A(_03185_ ), .ZN(_04889_ ) );
OR2_X1 _12211_ ( .A1(_03248_ ), .A2(_03251_ ), .ZN(_04890_ ) );
AOI21_X1 _12212_ ( .A(_04889_ ), .B1(_04890_ ), .B2(_03178_ ), .ZN(_04891_ ) );
XNOR2_X1 _12213_ ( .A(_03186_ ), .B(_03142_ ), .ZN(_04892_ ) );
OAI22_X1 _12214_ ( .A1(_04891_ ), .A2(_03195_ ), .B1(\u_exu.alu_p1[13] ), .B2(_04892_ ), .ZN(_04893_ ) );
AOI21_X1 _12215_ ( .A(_04888_ ), .B1(_04893_ ), .B2(_03194_ ), .ZN(_04894_ ) );
OR3_X1 _12216_ ( .A1(_04894_ ), .A2(_03149_ ), .A3(_03152_ ), .ZN(_04895_ ) );
OAI21_X1 _12217_ ( .A(_03149_ ), .B1(_04894_ ), .B2(_03152_ ), .ZN(_04896_ ) );
NAND3_X1 _12218_ ( .A1(_04895_ ), .A2(_04586_ ), .A3(_04896_ ), .ZN(_04897_ ) );
NAND3_X1 _12219_ ( .A1(_04530_ ), .A2(_04489_ ), .A3(_04502_ ), .ZN(_04898_ ) );
NOR2_X1 _12220_ ( .A1(_03418_ ), .A2(\u_exu.alu_ctrl[1] ), .ZN(_04899_ ) );
INV_X1 _12221_ ( .A(_04899_ ), .ZN(_04900_ ) );
NOR3_X1 _12222_ ( .A1(_04898_ ), .A2(fanout_net_19 ), .A3(_04900_ ), .ZN(_04901_ ) );
OR3_X1 _12223_ ( .A1(_04547_ ), .A2(_04482_ ), .A3(_04545_ ), .ZN(_04902_ ) );
OR3_X1 _12224_ ( .A1(_04511_ ), .A2(fanout_net_16 ), .A3(_04548_ ), .ZN(_04903_ ) );
NAND3_X1 _12225_ ( .A1(_04902_ ), .A2(_04903_ ), .A3(_04489_ ), .ZN(_04904_ ) );
NAND3_X1 _12226_ ( .A1(_04769_ ), .A2(_04770_ ), .A3(fanout_net_18 ), .ZN(_04905_ ) );
NAND2_X1 _12227_ ( .A1(_04904_ ), .A2(_04905_ ), .ZN(_04906_ ) );
AOI21_X1 _12228_ ( .A(fanout_net_18 ), .B1(_04772_ ), .B2(_04773_ ), .ZN(_04907_ ) );
AOI21_X1 _12229_ ( .A(_04907_ ), .B1(fanout_net_18 ), .B2(_04766_ ), .ZN(_04908_ ) );
MUX2_X1 _12230_ ( .A(_04906_ ), .B(_04908_ ), .S(fanout_net_19 ), .Z(_04909_ ) );
AOI21_X1 _12231_ ( .A(_04901_ ), .B1(_04909_ ), .B2(_04679_ ), .ZN(_04910_ ) );
AOI21_X1 _12232_ ( .A(_04571_ ), .B1(_04910_ ), .B2(_04677_ ), .ZN(_04911_ ) );
AND3_X1 _12233_ ( .A1(_04499_ ), .A2(_04521_ ), .A3(_04563_ ), .ZN(_04912_ ) );
NAND2_X1 _12234_ ( .A1(_03095_ ), .A2(_04574_ ), .ZN(_04913_ ) );
AOI21_X1 _12235_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[15] ), .B2(\u_exu.alu_p2[15] ), .ZN(_04914_ ) );
BUF_X4 _12236_ ( .A(_04565_ ), .Z(_04915_ ) );
OAI211_X1 _12237_ ( .A(_04915_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[15] ), .C2(\u_exu.alu_p2[15] ), .ZN(_04916_ ) );
OAI211_X1 _12238_ ( .A(_04913_ ), .B(_04577_ ), .C1(_04914_ ), .C2(_04916_ ), .ZN(_04917_ ) );
NOR3_X1 _12239_ ( .A1(_04911_ ), .A2(_04912_ ), .A3(_04917_ ), .ZN(_04918_ ) );
AOI211_X1 _12240_ ( .A(_04582_ ), .B(_04887_ ), .C1(_04897_ ), .C2(_04918_ ), .ZN(_00312_ ) );
AND4_X1 _12241_ ( .A1(_03179_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(fanout_net_20 ), .ZN(_04919_ ) );
AND3_X1 _12242_ ( .A1(_04893_ ), .A2(_04888_ ), .A3(_03194_ ), .ZN(_04920_ ) );
OR3_X1 _12243_ ( .A1(_04920_ ), .A2(_04894_ ), .A3(_04713_ ), .ZN(_04921_ ) );
NAND2_X1 _12244_ ( .A1(_03117_ ), .A2(_04639_ ), .ZN(_04922_ ) );
AOI21_X1 _12245_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[14] ), .B2(\u_exu.alu_p2[14] ), .ZN(_04923_ ) );
OAI211_X1 _12246_ ( .A(_04642_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[14] ), .C2(\u_exu.alu_p2[14] ), .ZN(_04924_ ) );
OAI211_X1 _12247_ ( .A(_04922_ ), .B(_03071_ ), .C1(_04923_ ), .C2(_04924_ ), .ZN(_04925_ ) );
AND3_X1 _12248_ ( .A1(_04598_ ), .A2(_04563_ ), .A3(_04607_ ), .ZN(_04926_ ) );
AND3_X1 _12249_ ( .A1(_04825_ ), .A2(_04826_ ), .A3(_03455_ ), .ZN(_04927_ ) );
AOI21_X1 _12250_ ( .A(_04927_ ), .B1(_04817_ ), .B2(fanout_net_18 ), .ZN(_04928_ ) );
AOI21_X1 _12251_ ( .A(_03456_ ), .B1(_04822_ ), .B2(_04823_ ), .ZN(_04929_ ) );
OR3_X1 _12252_ ( .A1(_03386_ ), .A2(_03387_ ), .A3(_04659_ ), .ZN(_04930_ ) );
OR3_X1 _12253_ ( .A1(_03437_ ), .A2(_03438_ ), .A3(fanout_net_16 ), .ZN(_04931_ ) );
AOI21_X1 _12254_ ( .A(fanout_net_18 ), .B1(_04930_ ), .B2(_04931_ ), .ZN(_04932_ ) );
NOR2_X1 _12255_ ( .A1(_04929_ ), .A2(_04932_ ), .ZN(_04933_ ) );
MUX2_X1 _12256_ ( .A(_04928_ ), .B(_04933_ ), .S(_04523_ ), .Z(_04934_ ) );
OR2_X1 _12257_ ( .A1(_04934_ ), .A2(\u_exu.alu_p2[4] ), .ZN(_04935_ ) );
INV_X1 _12258_ ( .A(_04615_ ), .ZN(_04936_ ) );
NOR3_X1 _12259_ ( .A1(_04612_ ), .A2(_04613_ ), .A3(_04936_ ), .ZN(_04937_ ) );
INV_X1 _12260_ ( .A(_04617_ ), .ZN(_04938_ ) );
AOI211_X1 _12261_ ( .A(_04571_ ), .B(_04937_ ), .C1(_04938_ ), .C2(_04899_ ), .ZN(_04939_ ) );
AOI211_X1 _12262_ ( .A(_04925_ ), .B(_04926_ ), .C1(_04935_ ), .C2(_04939_ ), .ZN(_04940_ ) );
AOI211_X1 _12263_ ( .A(_04582_ ), .B(_04919_ ), .C1(_04921_ ), .C2(_04940_ ), .ZN(_00313_ ) );
AND4_X1 _12264_ ( .A1(_03192_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(fanout_net_20 ), .ZN(_04941_ ) );
OR3_X1 _12265_ ( .A1(_04891_ ), .A2(_03195_ ), .A3(_03188_ ), .ZN(_04942_ ) );
OAI21_X1 _12266_ ( .A(_03188_ ), .B1(_04891_ ), .B2(_03195_ ), .ZN(_04943_ ) );
NAND3_X1 _12267_ ( .A1(_04942_ ), .A2(_04586_ ), .A3(_04943_ ), .ZN(_04944_ ) );
NOR2_X1 _12268_ ( .A1(_04663_ ), .A2(_04520_ ), .ZN(_04945_ ) );
NAND3_X1 _12269_ ( .A1(_04840_ ), .A2(_04841_ ), .A3(fanout_net_18 ), .ZN(_04946_ ) );
OR3_X1 _12270_ ( .A1(_04511_ ), .A2(_04659_ ), .A3(_04548_ ), .ZN(_04947_ ) );
OR3_X1 _12271_ ( .A1(_04514_ ), .A2(_04512_ ), .A3(fanout_net_16 ), .ZN(_04948_ ) );
NAND3_X1 _12272_ ( .A1(_04947_ ), .A2(_03456_ ), .A3(_04948_ ), .ZN(_04949_ ) );
AOI21_X1 _12273_ ( .A(fanout_net_19 ), .B1(_04946_ ), .B2(_04949_ ), .ZN(_04950_ ) );
OAI21_X1 _12274_ ( .A(_04679_ ), .B1(_04945_ ), .B2(_04950_ ), .ZN(_04951_ ) );
NOR2_X1 _12275_ ( .A1(_04613_ ), .A2(_03366_ ), .ZN(_04952_ ) );
OAI21_X1 _12276_ ( .A(_04952_ ), .B1(_04669_ ), .B2(fanout_net_19 ), .ZN(_04953_ ) );
OR3_X1 _12277_ ( .A1(_04673_ ), .A2(fanout_net_19 ), .A3(fanout_net_18 ), .ZN(_04954_ ) );
NAND2_X1 _12278_ ( .A1(_04954_ ), .A2(_03366_ ), .ZN(_04955_ ) );
NAND3_X1 _12279_ ( .A1(_04953_ ), .A2(\u_exu.alu_p2[4] ), .A3(_04955_ ), .ZN(_04956_ ) );
AOI21_X1 _12280_ ( .A(_04571_ ), .B1(_04951_ ), .B2(_04956_ ), .ZN(_04957_ ) );
OR2_X1 _12281_ ( .A1(_04705_ ), .A2(_04519_ ), .ZN(_04958_ ) );
NAND3_X1 _12282_ ( .A1(_04683_ ), .A2(_04687_ ), .A3(_04523_ ), .ZN(_04959_ ) );
AND3_X1 _12283_ ( .A1(_04958_ ), .A2(_04563_ ), .A3(_04959_ ), .ZN(_04960_ ) );
OAI211_X1 _12284_ ( .A(_04642_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[13] ), .C2(\u_exu.alu_p2[13] ), .ZN(_04961_ ) );
INV_X1 _12285_ ( .A(\u_exu.alu_ctrl[0] ), .ZN(_04962_ ) );
NAND2_X1 _12286_ ( .A1(\u_exu.alu_p1[13] ), .A2(\u_exu.alu_p2[13] ), .ZN(_04963_ ) );
AOI21_X1 _12287_ ( .A(_04961_ ), .B1(_04962_ ), .B2(_04963_ ), .ZN(_04964_ ) );
NAND2_X1 _12288_ ( .A1(_03115_ ), .A2(_04639_ ), .ZN(_04965_ ) );
NAND2_X1 _12289_ ( .A1(_04965_ ), .A2(_03071_ ), .ZN(_04966_ ) );
NOR4_X1 _12290_ ( .A1(_04957_ ), .A2(_04960_ ), .A3(_04964_ ), .A4(_04966_ ), .ZN(_04967_ ) );
AOI211_X1 _12291_ ( .A(_04582_ ), .B(_04941_ ), .C1(_04944_ ), .C2(_04967_ ), .ZN(_00314_ ) );
AND3_X1 _12292_ ( .A1(_04890_ ), .A2(_04889_ ), .A3(_03178_ ), .ZN(_04968_ ) );
OR3_X1 _12293_ ( .A1(_04968_ ), .A2(_04891_ ), .A3(_04712_ ), .ZN(_04969_ ) );
OR2_X1 _12294_ ( .A1(_04752_ ), .A2(_03453_ ), .ZN(_04970_ ) );
NAND2_X1 _12295_ ( .A1(_04735_ ), .A2(_04518_ ), .ZN(_04971_ ) );
AND3_X1 _12296_ ( .A1(_04970_ ), .A2(_04562_ ), .A3(_04971_ ), .ZN(_04972_ ) );
NOR3_X1 _12297_ ( .A1(_04721_ ), .A2(_04722_ ), .A3(_03453_ ), .ZN(_04973_ ) );
AOI21_X1 _12298_ ( .A(_03456_ ), .B1(_03385_ ), .B2(_03388_ ), .ZN(_04974_ ) );
AND3_X1 _12299_ ( .A1(_03436_ ), .A2(_03439_ ), .A3(_03455_ ), .ZN(_04975_ ) );
NOR2_X1 _12300_ ( .A1(_04974_ ), .A2(_04975_ ), .ZN(_04976_ ) );
AOI21_X1 _12301_ ( .A(_04973_ ), .B1(_03454_ ), .B2(_04976_ ), .ZN(_04977_ ) );
AOI21_X1 _12302_ ( .A(_03381_ ), .B1(_04977_ ), .B2(_04679_ ), .ZN(_04978_ ) );
INV_X1 _12303_ ( .A(_04952_ ), .ZN(_04979_ ) );
AOI21_X1 _12304_ ( .A(_04979_ ), .B1(_04719_ ), .B2(_03454_ ), .ZN(_04980_ ) );
NOR3_X1 _12305_ ( .A1(_03414_ ), .A2(\u_exu.alu_p2[3] ), .A3(\u_exu.alu_p2[2] ), .ZN(_04981_ ) );
NOR2_X1 _12306_ ( .A1(_04981_ ), .A2(\u_exu.alu_ctrl[1] ), .ZN(_04982_ ) );
OAI21_X1 _12307_ ( .A(\u_exu.alu_p2[4] ), .B1(_04980_ ), .B2(_04982_ ), .ZN(_04983_ ) );
AOI221_X4 _12308_ ( .A(_04972_ ), .B1(_03092_ ), .B2(_04573_ ), .C1(_04978_ ), .C2(_04983_ ), .ZN(_04984_ ) );
AOI21_X1 _12309_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[12] ), .B2(\u_exu.alu_p2[12] ), .ZN(_04985_ ) );
OAI211_X1 _12310_ ( .A(_04915_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[12] ), .C2(\u_exu.alu_p2[12] ), .ZN(_04986_ ) );
OAI211_X1 _12311_ ( .A(_04969_ ), .B(_04984_ ), .C1(_04985_ ), .C2(_04986_ ), .ZN(_04987_ ) );
MUX2_X1 _12312_ ( .A(\u_exu.alu_p1[12] ), .B(_04987_ ), .S(_04577_ ), .Z(_04988_ ) );
AND2_X1 _12313_ ( .A1(_04988_ ), .A2(_04580_ ), .ZN(_00315_ ) );
NOR2_X1 _12314_ ( .A1(_03350_ ), .A2(\u_exu.alu_p1[28] ), .ZN(_04989_ ) );
NOR3_X1 _12315_ ( .A1(_03343_ ), .A2(_03354_ ), .A3(_04989_ ), .ZN(_04990_ ) );
OR3_X1 _12316_ ( .A1(_04990_ ), .A2(_03348_ ), .A3(_03354_ ), .ZN(_04991_ ) );
OAI21_X1 _12317_ ( .A(_03348_ ), .B1(_04990_ ), .B2(_03354_ ), .ZN(_04992_ ) );
NAND3_X1 _12318_ ( .A1(_04991_ ), .A2(_04586_ ), .A3(_04992_ ), .ZN(_04993_ ) );
NOR4_X1 _12319_ ( .A1(_03129_ ), .A2(_03379_ ), .A3(_03373_ ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_04994_ ) );
OAI21_X1 _12320_ ( .A(_04994_ ), .B1(\u_exu.alu_ctrl[0] ), .B2(_03128_ ), .ZN(_04995_ ) );
NAND3_X1 _12321_ ( .A1(_03130_ ), .A2(fanout_net_20 ), .A3(_03083_ ), .ZN(_04996_ ) );
MUX2_X1 _12322_ ( .A(\u_exu.alu_p1[31] ), .B(_04953_ ), .S(_03418_ ), .Z(_04997_ ) );
AND2_X1 _12323_ ( .A1(_03380_ ), .A2(_04900_ ), .ZN(_04998_ ) );
NAND3_X1 _12324_ ( .A1(_04997_ ), .A2(_04955_ ), .A3(_04998_ ), .ZN(_04999_ ) );
NAND3_X1 _12325_ ( .A1(_04958_ ), .A2(_04501_ ), .A3(_04959_ ), .ZN(_05000_ ) );
NAND3_X1 _12326_ ( .A1(_04556_ ), .A2(fanout_net_16 ), .A3(_04558_ ), .ZN(_05001_ ) );
NAND3_X1 _12327_ ( .A1(_04538_ ), .A2(_04528_ ), .A3(_04540_ ), .ZN(_05002_ ) );
AOI21_X1 _12328_ ( .A(_03457_ ), .B1(_05001_ ), .B2(_05002_ ), .ZN(_05003_ ) );
NOR2_X1 _12329_ ( .A1(_04655_ ), .A2(_04534_ ), .ZN(_05004_ ) );
MUX2_X1 _12330_ ( .A(_05004_ ), .B(_04527_ ), .S(_04528_ ), .Z(_05005_ ) );
AOI211_X1 _12331_ ( .A(\u_exu.alu_p2[3] ), .B(_05003_ ), .C1(_04498_ ), .C2(_05005_ ), .ZN(_05006_ ) );
AOI21_X1 _12332_ ( .A(_04523_ ), .B1(_04694_ ), .B2(_04697_ ), .ZN(_05007_ ) );
OAI21_X1 _12333_ ( .A(_04637_ ), .B1(_05006_ ), .B2(_05007_ ), .ZN(_05008_ ) );
AND3_X1 _12334_ ( .A1(_04999_ ), .A2(_05000_ ), .A3(_05008_ ), .ZN(_05009_ ) );
NAND4_X1 _12335_ ( .A1(_04993_ ), .A2(_04995_ ), .A3(_04996_ ), .A4(_05009_ ), .ZN(_05010_ ) );
MUX2_X1 _12336_ ( .A(\u_exu.alu_p1[29] ), .B(_05010_ ), .S(_04578_ ), .Z(_05011_ ) );
AND2_X1 _12337_ ( .A1(_05011_ ), .A2(_04580_ ), .ZN(_00316_ ) );
NOR4_X1 _12338_ ( .A1(_03379_ ), .A2(\u_exu.alu_p1[11] ), .A3(\u_exu.alu_ctrl[5] ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_05012_ ) );
INV_X1 _12339_ ( .A(_03176_ ), .ZN(_05013_ ) );
INV_X1 _12340_ ( .A(_03250_ ), .ZN(_05014_ ) );
NOR2_X1 _12341_ ( .A1(_03248_ ), .A2(_05014_ ), .ZN(_05015_ ) );
AND2_X1 _12342_ ( .A1(_05015_ ), .A2(_03167_ ), .ZN(_05016_ ) );
INV_X1 _12343_ ( .A(_05016_ ), .ZN(_05017_ ) );
AOI21_X1 _12344_ ( .A(_05013_ ), .B1(_05017_ ), .B2(_03173_ ), .ZN(_05018_ ) );
OR3_X1 _12345_ ( .A1(_05018_ ), .A2(_03158_ ), .A3(_03161_ ), .ZN(_05019_ ) );
OAI21_X1 _12346_ ( .A(_03158_ ), .B1(_05018_ ), .B2(_03161_ ), .ZN(_05020_ ) );
NAND3_X1 _12347_ ( .A1(_05019_ ), .A2(_04586_ ), .A3(_05020_ ), .ZN(_05021_ ) );
NAND3_X1 _12348_ ( .A1(_04902_ ), .A2(_04903_ ), .A3(\u_exu.alu_p2[2] ), .ZN(_05022_ ) );
OR3_X1 _12349_ ( .A1(_04503_ ), .A2(fanout_net_16 ), .A3(_04515_ ), .ZN(_05023_ ) );
OR3_X1 _12350_ ( .A1(_04514_ ), .A2(_04512_ ), .A3(_04482_ ), .ZN(_05024_ ) );
NAND3_X1 _12351_ ( .A1(_05023_ ), .A2(_03455_ ), .A3(_05024_ ), .ZN(_05025_ ) );
AND2_X1 _12352_ ( .A1(_05022_ ), .A2(_05025_ ), .ZN(_05026_ ) );
AND2_X1 _12353_ ( .A1(_04771_ ), .A2(_04774_ ), .ZN(_05027_ ) );
MUX2_X1 _12354_ ( .A(_05026_ ), .B(_05027_ ), .S(\u_exu.alu_p2[3] ), .Z(_05028_ ) );
AOI21_X1 _12355_ ( .A(\u_exu.alu_p2[3] ), .B1(_04767_ ), .B2(_04718_ ), .ZN(_05029_ ) );
NOR2_X1 _12356_ ( .A1(_05029_ ), .A2(_04979_ ), .ZN(_05030_ ) );
MUX2_X1 _12357_ ( .A(_05028_ ), .B(_05030_ ), .S(\u_exu.alu_p2[4] ), .Z(_05031_ ) );
INV_X1 _12358_ ( .A(_04998_ ), .ZN(_05032_ ) );
NAND3_X1 _12359_ ( .A1(_04778_ ), .A2(_04524_ ), .A3(_04717_ ), .ZN(_05033_ ) );
AOI21_X1 _12360_ ( .A(_05031_ ), .B1(_05032_ ), .B2(_05033_ ), .ZN(_05034_ ) );
OAI21_X1 _12361_ ( .A(\u_exu.alu_p2[3] ), .B1(_04497_ ), .B2(\u_exu.alu_p2[2] ), .ZN(_05035_ ) );
NAND3_X1 _12362_ ( .A1(_04783_ ), .A2(_04784_ ), .A3(_04519_ ), .ZN(_05036_ ) );
AND3_X1 _12363_ ( .A1(_05035_ ), .A2(_05036_ ), .A3(_04563_ ), .ZN(_05037_ ) );
NAND2_X1 _12364_ ( .A1(_04574_ ), .A2(_03118_ ), .ZN(_05038_ ) );
AOI21_X1 _12365_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[11] ), .B2(\u_exu.alu_p2[11] ), .ZN(_05039_ ) );
OAI211_X1 _12366_ ( .A(_04915_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[11] ), .C2(\u_exu.alu_p2[11] ), .ZN(_05040_ ) );
OAI211_X1 _12367_ ( .A(_05038_ ), .B(_04577_ ), .C1(_05039_ ), .C2(_05040_ ), .ZN(_05041_ ) );
NOR3_X1 _12368_ ( .A1(_05034_ ), .A2(_05037_ ), .A3(_05041_ ), .ZN(_05042_ ) );
AOI211_X1 _12369_ ( .A(_04582_ ), .B(_05012_ ), .C1(_05021_ ), .C2(_05042_ ), .ZN(_00317_ ) );
AND4_X1 _12370_ ( .A1(_03175_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(fanout_net_20 ), .ZN(_05043_ ) );
AOI211_X1 _12371_ ( .A(_03176_ ), .B(_03174_ ), .C1(_05015_ ), .C2(_03167_ ), .ZN(_05044_ ) );
OR3_X1 _12372_ ( .A1(_05018_ ), .A2(_04713_ ), .A3(_05044_ ), .ZN(_05045_ ) );
NOR3_X1 _12373_ ( .A1(_04824_ ), .A2(_04827_ ), .A3(_04599_ ), .ZN(_05046_ ) );
OR3_X1 _12374_ ( .A1(_03434_ ), .A2(_03435_ ), .A3(_04482_ ), .ZN(_05047_ ) );
OR3_X1 _12375_ ( .A1(_03442_ ), .A2(_03443_ ), .A3(fanout_net_16 ), .ZN(_05048_ ) );
NAND3_X1 _12376_ ( .A1(_05047_ ), .A2(_05048_ ), .A3(_03457_ ), .ZN(_05049_ ) );
NAND3_X1 _12377_ ( .A1(_04930_ ), .A2(_04931_ ), .A3(\u_exu.alu_p2[2] ), .ZN(_05050_ ) );
NAND2_X1 _12378_ ( .A1(_05049_ ), .A2(_05050_ ), .ZN(_05051_ ) );
AOI211_X1 _12379_ ( .A(\u_exu.alu_p2[4] ), .B(_05046_ ), .C1(_04600_ ), .C2(_05051_ ), .ZN(_05052_ ) );
AND2_X1 _12380_ ( .A1(_04818_ ), .A2(_03454_ ), .ZN(_05053_ ) );
AOI21_X1 _12381_ ( .A(_04998_ ), .B1(_05053_ ), .B2(_03380_ ), .ZN(_05054_ ) );
OR2_X1 _12382_ ( .A1(_05052_ ), .A2(_05054_ ), .ZN(_05055_ ) );
OAI21_X1 _12383_ ( .A(_03453_ ), .B1(_04818_ ), .B2(_04819_ ), .ZN(_05056_ ) );
AND2_X1 _12384_ ( .A1(_05056_ ), .A2(_04952_ ), .ZN(_05057_ ) );
AOI21_X1 _12385_ ( .A(_05055_ ), .B1(\u_exu.alu_p2[4] ), .B2(_05057_ ), .ZN(_05058_ ) );
OAI21_X1 _12386_ ( .A(_04599_ ), .B1(_04800_ ), .B2(_04801_ ), .ZN(_05059_ ) );
OAI21_X1 _12387_ ( .A(\u_exu.alu_p2[3] ), .B1(_04596_ ), .B2(\u_exu.alu_p2[2] ), .ZN(_05060_ ) );
AND3_X1 _12388_ ( .A1(_05059_ ), .A2(_04563_ ), .A3(_05060_ ), .ZN(_05061_ ) );
NAND2_X1 _12389_ ( .A1(_03093_ ), .A2(_04574_ ), .ZN(_05062_ ) );
AOI21_X1 _12390_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[10] ), .B2(\u_exu.alu_p2[10] ), .ZN(_05063_ ) );
OAI211_X1 _12391_ ( .A(_04915_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[10] ), .C2(\u_exu.alu_p2[10] ), .ZN(_05064_ ) );
OAI211_X1 _12392_ ( .A(_05062_ ), .B(_03071_ ), .C1(_05063_ ), .C2(_05064_ ), .ZN(_05065_ ) );
NOR3_X1 _12393_ ( .A1(_05058_ ), .A2(_05061_ ), .A3(_05065_ ), .ZN(_05066_ ) );
AOI211_X1 _12394_ ( .A(_04451_ ), .B(_05043_ ), .C1(_05045_ ), .C2(_05066_ ), .ZN(_00318_ ) );
NOR4_X1 _12395_ ( .A1(_03379_ ), .A2(\u_exu.alu_p1[9] ), .A3(\u_exu.alu_ctrl[5] ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_05067_ ) );
OR3_X1 _12396_ ( .A1(_05015_ ), .A2(_03167_ ), .A3(_03170_ ), .ZN(_05068_ ) );
OAI21_X1 _12397_ ( .A(_03167_ ), .B1(_05015_ ), .B2(_03170_ ), .ZN(_05069_ ) );
NAND3_X1 _12398_ ( .A1(_05068_ ), .A2(_04586_ ), .A3(_05069_ ), .ZN(_05070_ ) );
NOR2_X1 _12399_ ( .A1(_04848_ ), .A2(\u_exu.alu_p2[3] ), .ZN(_05071_ ) );
NOR2_X1 _12400_ ( .A1(_04838_ ), .A2(\u_exu.alu_p2[3] ), .ZN(_05072_ ) );
OAI22_X1 _12401_ ( .A1(_05071_ ), .A2(_04979_ ), .B1(\u_exu.alu_ctrl[1] ), .B2(_05072_ ), .ZN(_05073_ ) );
AND2_X1 _12402_ ( .A1(_05073_ ), .A2(\u_exu.alu_p2[4] ), .ZN(_05074_ ) );
OR3_X1 _12403_ ( .A1(_04503_ ), .A2(_04659_ ), .A3(_04515_ ), .ZN(_05075_ ) );
OR3_X1 _12404_ ( .A1(_04506_ ), .A2(fanout_net_16 ), .A3(_04504_ ), .ZN(_05076_ ) );
AOI21_X1 _12405_ ( .A(\u_exu.alu_p2[2] ), .B1(_05075_ ), .B2(_05076_ ), .ZN(_05077_ ) );
AOI21_X1 _12406_ ( .A(_04490_ ), .B1(_04947_ ), .B2(_04948_ ), .ZN(_05078_ ) );
OAI21_X1 _12407_ ( .A(_04600_ ), .B1(_05077_ ), .B2(_05078_ ), .ZN(_05079_ ) );
NAND3_X1 _12408_ ( .A1(_04842_ ), .A2(_04843_ ), .A3(\u_exu.alu_p2[3] ), .ZN(_05080_ ) );
AOI21_X1 _12409_ ( .A(\u_exu.alu_p2[4] ), .B1(_05079_ ), .B2(_05080_ ), .ZN(_05081_ ) );
OR3_X1 _12410_ ( .A1(_05074_ ), .A2(_04571_ ), .A3(_05081_ ), .ZN(_05082_ ) );
OAI211_X1 _12411_ ( .A(_04642_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p2[9] ), .C2(\u_exu.alu_p1[9] ), .ZN(_05083_ ) );
NAND2_X1 _12412_ ( .A1(\u_exu.alu_p2[9] ), .A2(\u_exu.alu_p1[9] ), .ZN(_05084_ ) );
AOI21_X1 _12413_ ( .A(_05083_ ), .B1(_04962_ ), .B2(_05084_ ), .ZN(_05085_ ) );
NAND2_X1 _12414_ ( .A1(_04858_ ), .A2(_04519_ ), .ZN(_05086_ ) );
OR2_X1 _12415_ ( .A1(_04860_ ), .A2(_03454_ ), .ZN(_05087_ ) );
AND3_X1 _12416_ ( .A1(_05086_ ), .A2(_04637_ ), .A3(_05087_ ), .ZN(_05088_ ) );
AOI211_X1 _12417_ ( .A(_05085_ ), .B(_05088_ ), .C1(_03094_ ), .C2(_04574_ ), .ZN(_05089_ ) );
AND3_X1 _12418_ ( .A1(_05082_ ), .A2(_04577_ ), .A3(_05089_ ), .ZN(_05090_ ) );
AOI211_X1 _12419_ ( .A(_04451_ ), .B(_05067_ ), .C1(_05070_ ), .C2(_05090_ ), .ZN(_00319_ ) );
OAI21_X1 _12420_ ( .A(_04478_ ), .B1(_03248_ ), .B2(_05014_ ), .ZN(_05091_ ) );
AOI21_X1 _12421_ ( .A(_05091_ ), .B1(_03248_ ), .B2(_05014_ ), .ZN(_05092_ ) );
OAI211_X1 _12422_ ( .A(_04565_ ), .B(fanout_net_20 ), .C1(\u_exu.alu_p1[8] ), .C2(\u_exu.alu_p2[8] ), .ZN(_05093_ ) );
NAND2_X1 _12423_ ( .A1(\u_exu.alu_p1[8] ), .A2(\u_exu.alu_p2[8] ), .ZN(_05094_ ) );
AOI21_X1 _12424_ ( .A(_05093_ ), .B1(_04962_ ), .B2(_05094_ ), .ZN(_05095_ ) );
AND2_X1 _12425_ ( .A1(_03116_ ), .A2(_04639_ ), .ZN(_05096_ ) );
AND2_X1 _12426_ ( .A1(_03415_ ), .A2(_04518_ ), .ZN(_05097_ ) );
INV_X1 _12427_ ( .A(_05097_ ), .ZN(_05098_ ) );
AOI21_X1 _12428_ ( .A(_03418_ ), .B1(_04613_ ), .B2(\u_exu.alu_ctrl[1] ), .ZN(_05099_ ) );
AOI21_X1 _12429_ ( .A(_03381_ ), .B1(_05098_ ), .B2(_05099_ ), .ZN(_05100_ ) );
NAND2_X1 _12430_ ( .A1(_03441_ ), .A2(_03448_ ), .ZN(_05101_ ) );
MUX2_X1 _12431_ ( .A(_05101_ ), .B(_03398_ ), .S(\u_exu.alu_p2[3] ), .Z(_05102_ ) );
OAI21_X1 _12432_ ( .A(_05100_ ), .B1(\u_exu.alu_p2[4] ), .B2(_05102_ ), .ZN(_05103_ ) );
NAND3_X1 _12433_ ( .A1(_04874_ ), .A2(_04875_ ), .A3(_04599_ ), .ZN(_05104_ ) );
NAND4_X1 _12434_ ( .A1(_03420_ ), .A2(\u_exu.alu_p2[3] ), .A3(_03457_ ), .A4(_04528_ ), .ZN(_05105_ ) );
AOI21_X1 _12435_ ( .A(\u_exu.alu_p2[4] ), .B1(_05104_ ), .B2(_05105_ ), .ZN(_05106_ ) );
NAND2_X1 _12436_ ( .A1(_05106_ ), .A2(_03378_ ), .ZN(_05107_ ) );
NAND2_X1 _12437_ ( .A1(_05103_ ), .A2(_05107_ ), .ZN(_05108_ ) );
NOR4_X1 _12438_ ( .A1(_05092_ ), .A2(_05095_ ), .A3(_05096_ ), .A4(_05108_ ), .ZN(_05109_ ) );
MUX2_X1 _12439_ ( .A(_03249_ ), .B(_05109_ ), .S(_04577_ ), .Z(_05110_ ) );
OR2_X1 _12440_ ( .A1(_05110_ ), .A2(_01075_ ), .ZN(_05111_ ) );
INV_X1 _12441_ ( .A(_05111_ ), .ZN(_00320_ ) );
AND4_X1 _12442_ ( .A1(\u_exu.alu_p1[7] ), .A2(_04583_ ), .A3(_04584_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05112_ ) );
AOI21_X1 _12443_ ( .A(_03219_ ), .B1(_03235_ ), .B2(_03239_ ), .ZN(_05113_ ) );
INV_X1 _12444_ ( .A(_03246_ ), .ZN(_05114_ ) );
OAI21_X1 _12445_ ( .A(_03204_ ), .B1(_05113_ ), .B2(_05114_ ), .ZN(_05115_ ) );
NAND2_X1 _12446_ ( .A1(_03202_ ), .A2(\u_exu.alu_p1[6] ), .ZN(_05116_ ) );
AND3_X1 _12447_ ( .A1(_05115_ ), .A2(_03209_ ), .A3(_05116_ ), .ZN(_05117_ ) );
AOI21_X1 _12448_ ( .A(_03209_ ), .B1(_05115_ ), .B2(_05116_ ), .ZN(_05118_ ) );
OAI21_X1 _12449_ ( .A(_04478_ ), .B1(_05117_ ), .B2(_05118_ ), .ZN(_05119_ ) );
NOR3_X1 _12450_ ( .A1(_04898_ ), .A2(\u_exu.alu_ctrl[1] ), .A3(_04518_ ), .ZN(_05120_ ) );
AOI21_X1 _12451_ ( .A(_05120_ ), .B1(_04908_ ), .B2(_04519_ ), .ZN(_05121_ ) );
AOI21_X1 _12452_ ( .A(_03381_ ), .B1(_05121_ ), .B2(_05099_ ), .ZN(_05122_ ) );
NAND3_X1 _12453_ ( .A1(_05023_ ), .A2(\u_exu.alu_p2[2] ), .A3(_05024_ ), .ZN(_05123_ ) );
OAI21_X1 _12454_ ( .A(_04482_ ), .B1(_04486_ ), .B2(_04507_ ), .ZN(_05124_ ) );
OAI21_X1 _12455_ ( .A(fanout_net_16 ), .B1(_04506_ ), .B2(_04504_ ), .ZN(_05125_ ) );
AND2_X1 _12456_ ( .A1(_05124_ ), .A2(_05125_ ), .ZN(_05126_ ) );
OAI21_X1 _12457_ ( .A(_05123_ ), .B1(_05126_ ), .B2(\u_exu.alu_p2[2] ), .ZN(_05127_ ) );
MUX2_X1 _12458_ ( .A(_04906_ ), .B(_05127_ ), .S(_04599_ ), .Z(_05128_ ) );
OAI21_X1 _12459_ ( .A(_05122_ ), .B1(\u_exu.alu_p2[4] ), .B2(_05128_ ), .ZN(_05129_ ) );
OAI21_X1 _12460_ ( .A(_04491_ ), .B1(_04497_ ), .B2(_04498_ ), .ZN(_05130_ ) );
NAND3_X1 _12461_ ( .A1(_05130_ ), .A2(_04520_ ), .A3(_04637_ ), .ZN(_05131_ ) );
NAND2_X1 _12462_ ( .A1(_04639_ ), .A2(_03087_ ), .ZN(_05132_ ) );
AND3_X1 _12463_ ( .A1(_05129_ ), .A2(_05131_ ), .A3(_05132_ ), .ZN(_05133_ ) );
AOI21_X1 _12464_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[7] ), .B2(\u_exu.alu_p2[7] ), .ZN(_05134_ ) );
OAI211_X1 _12465_ ( .A(_04915_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[7] ), .C2(\u_exu.alu_p2[7] ), .ZN(_05135_ ) );
OAI211_X1 _12466_ ( .A(_05119_ ), .B(_05133_ ), .C1(_05134_ ), .C2(_05135_ ), .ZN(_05136_ ) );
AOI21_X1 _12467_ ( .A(_05112_ ), .B1(_05136_ ), .B2(_04578_ ), .ZN(_05137_ ) );
NOR2_X1 _12468_ ( .A1(_05137_ ), .A2(_04475_ ), .ZN(_00321_ ) );
OR3_X1 _12469_ ( .A1(_05113_ ), .A2(_03204_ ), .A3(_05114_ ), .ZN(_05138_ ) );
NAND3_X1 _12470_ ( .A1(_05138_ ), .A2(_04478_ ), .A3(_05115_ ), .ZN(_05139_ ) );
AND3_X1 _12471_ ( .A1(_04597_ ), .A2(_04599_ ), .A3(_04562_ ), .ZN(_05140_ ) );
AND2_X1 _12472_ ( .A1(_04928_ ), .A2(_03453_ ), .ZN(_05141_ ) );
NOR4_X1 _12473_ ( .A1(_03411_ ), .A2(_03453_ ), .A3(\u_exu.alu_p2[2] ), .A4(fanout_net_16 ), .ZN(_05142_ ) );
OAI21_X1 _12474_ ( .A(_04899_ ), .B1(_05141_ ), .B2(_05142_ ), .ZN(_05143_ ) );
AOI21_X1 _12475_ ( .A(_03453_ ), .B1(_04610_ ), .B2(_04611_ ), .ZN(_05144_ ) );
OAI21_X1 _12476_ ( .A(_04615_ ), .B1(_05141_ ), .B2(_05144_ ), .ZN(_05145_ ) );
OR3_X1 _12477_ ( .A1(_03445_ ), .A2(_03446_ ), .A3(_04659_ ), .ZN(_05146_ ) );
OR3_X1 _12478_ ( .A1(_03425_ ), .A2(_03426_ ), .A3(fanout_net_16 ), .ZN(_05147_ ) );
AOI21_X1 _12479_ ( .A(\u_exu.alu_p2[2] ), .B1(_05146_ ), .B2(_05147_ ), .ZN(_05148_ ) );
AOI21_X1 _12480_ ( .A(_03456_ ), .B1(_05047_ ), .B2(_05048_ ), .ZN(_05149_ ) );
OAI21_X1 _12481_ ( .A(_04518_ ), .B1(_05148_ ), .B2(_05149_ ), .ZN(_05150_ ) );
OAI21_X1 _12482_ ( .A(_05150_ ), .B1(_04933_ ), .B2(_03454_ ), .ZN(_05151_ ) );
OAI211_X1 _12483_ ( .A(_05143_ ), .B(_05145_ ), .C1(\u_exu.alu_p2[4] ), .C2(_05151_ ), .ZN(_05152_ ) );
AOI221_X4 _12484_ ( .A(_05140_ ), .B1(_03111_ ), .B2(_04573_ ), .C1(_05152_ ), .C2(_04717_ ), .ZN(_05153_ ) );
AOI21_X1 _12485_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[6] ), .B2(\u_exu.alu_p2[6] ), .ZN(_05154_ ) );
OAI211_X1 _12486_ ( .A(_04915_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[6] ), .C2(\u_exu.alu_p2[6] ), .ZN(_05155_ ) );
OAI211_X1 _12487_ ( .A(_05139_ ), .B(_05153_ ), .C1(_05154_ ), .C2(_05155_ ), .ZN(_05156_ ) );
MUX2_X1 _12488_ ( .A(\u_exu.alu_p1[6] ), .B(_05156_ ), .S(_04578_ ), .Z(_05157_ ) );
AND2_X1 _12489_ ( .A1(_05157_ ), .A2(_04580_ ), .ZN(_00322_ ) );
INV_X1 _12490_ ( .A(_03214_ ), .ZN(_05158_ ) );
AOI21_X1 _12491_ ( .A(_05158_ ), .B1(_03235_ ), .B2(_03239_ ), .ZN(_05159_ ) );
OR3_X1 _12492_ ( .A1(_05159_ ), .A2(_03217_ ), .A3(_03245_ ), .ZN(_05160_ ) );
OAI21_X1 _12493_ ( .A(_03217_ ), .B1(_05159_ ), .B2(_03245_ ), .ZN(_05161_ ) );
NAND3_X1 _12494_ ( .A1(_05160_ ), .A2(_04478_ ), .A3(_05161_ ), .ZN(_05162_ ) );
AND3_X1 _12495_ ( .A1(_04705_ ), .A2(_04599_ ), .A3(_04562_ ), .ZN(_05163_ ) );
OAI21_X1 _12496_ ( .A(_04615_ ), .B1(_04664_ ), .B2(_04670_ ), .ZN(_05164_ ) );
OAI21_X1 _12497_ ( .A(_04899_ ), .B1(_04664_ ), .B2(_04674_ ), .ZN(_05165_ ) );
NAND3_X1 _12498_ ( .A1(_05075_ ), .A2(_05076_ ), .A3(\u_exu.alu_p2[2] ), .ZN(_05166_ ) );
OAI21_X1 _12499_ ( .A(_04483_ ), .B1(_04481_ ), .B2(_04487_ ), .ZN(_05167_ ) );
OAI21_X1 _12500_ ( .A(fanout_net_16 ), .B1(_04486_ ), .B2(_04507_ ), .ZN(_05168_ ) );
AND2_X1 _12501_ ( .A1(_05167_ ), .A2(_05168_ ), .ZN(_05169_ ) );
OAI211_X1 _12502_ ( .A(_05166_ ), .B(_04518_ ), .C1(\u_exu.alu_p2[2] ), .C2(_05169_ ), .ZN(_05170_ ) );
NAND3_X1 _12503_ ( .A1(_04946_ ), .A2(_04949_ ), .A3(\u_exu.alu_p2[3] ), .ZN(_05171_ ) );
NAND2_X1 _12504_ ( .A1(_05170_ ), .A2(_05171_ ), .ZN(_05172_ ) );
OAI211_X1 _12505_ ( .A(_05164_ ), .B(_05165_ ), .C1(\u_exu.alu_p2[4] ), .C2(_05172_ ), .ZN(_05173_ ) );
AOI221_X4 _12506_ ( .A(_05163_ ), .B1(_03113_ ), .B2(_04573_ ), .C1(_05173_ ), .C2(_03380_ ), .ZN(_05174_ ) );
AOI21_X1 _12507_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[5] ), .B2(\u_exu.alu_p2[5] ), .ZN(_05175_ ) );
OAI211_X1 _12508_ ( .A(_04915_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[5] ), .C2(\u_exu.alu_p2[5] ), .ZN(_05176_ ) );
OAI211_X1 _12509_ ( .A(_05162_ ), .B(_05174_ ), .C1(_05175_ ), .C2(_05176_ ), .ZN(_05177_ ) );
MUX2_X1 _12510_ ( .A(\u_exu.alu_p1[5] ), .B(_05177_ ), .S(_04577_ ), .Z(_05178_ ) );
AND2_X1 _12511_ ( .A1(_05178_ ), .A2(_04580_ ), .ZN(_00323_ ) );
AND4_X1 _12512_ ( .A1(_03213_ ), .A2(_03373_ ), .A3(_03077_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05179_ ) );
OAI21_X1 _12513_ ( .A(_04615_ ), .B1(_04720_ ), .B2(_04723_ ), .ZN(_05180_ ) );
OAI21_X1 _12514_ ( .A(_04899_ ), .B1(_04723_ ), .B2(_04725_ ), .ZN(_05181_ ) );
NAND3_X1 _12515_ ( .A1(_03444_ ), .A2(_03447_ ), .A3(\u_exu.alu_p2[2] ), .ZN(_05182_ ) );
OAI211_X1 _12516_ ( .A(_05182_ ), .B(_03454_ ), .C1(_03431_ ), .C2(\u_exu.alu_p2[2] ), .ZN(_05183_ ) );
OAI21_X1 _12517_ ( .A(_05183_ ), .B1(_04976_ ), .B2(_04519_ ), .ZN(_05184_ ) );
OAI211_X1 _12518_ ( .A(_05180_ ), .B(_05181_ ), .C1(\u_exu.alu_p2[4] ), .C2(_05184_ ), .ZN(_05185_ ) );
NAND2_X1 _12519_ ( .A1(_05185_ ), .A2(_04717_ ), .ZN(_05186_ ) );
NAND3_X1 _12520_ ( .A1(_04752_ ), .A2(_04520_ ), .A3(_04637_ ), .ZN(_05187_ ) );
INV_X1 _12521_ ( .A(_03460_ ), .ZN(_05188_ ) );
AOI21_X1 _12522_ ( .A(_05188_ ), .B1(_04962_ ), .B2(_03213_ ), .ZN(_05189_ ) );
AND2_X1 _12523_ ( .A1(\u_exu.alu_ctrl[0] ), .A2(\u_exu.alu_p1[4] ), .ZN(_05190_ ) );
OAI21_X1 _12524_ ( .A(_05189_ ), .B1(\u_exu.alu_p2[4] ), .B2(_05190_ ), .ZN(_05191_ ) );
AOI21_X1 _12525_ ( .A(_03070_ ), .B1(_03085_ ), .B2(_04639_ ), .ZN(_05192_ ) );
AND4_X1 _12526_ ( .A1(_05186_ ), .A2(_05187_ ), .A3(_05191_ ), .A4(_05192_ ), .ZN(_05193_ ) );
AND3_X1 _12527_ ( .A1(_03235_ ), .A2(_03239_ ), .A3(_05158_ ), .ZN(_05194_ ) );
OR3_X1 _12528_ ( .A1(_05194_ ), .A2(_05159_ ), .A3(_04713_ ), .ZN(_05195_ ) );
AOI211_X1 _12529_ ( .A(_04451_ ), .B(_05179_ ), .C1(_05193_ ), .C2(_05195_ ), .ZN(_00324_ ) );
AND3_X1 _12530_ ( .A1(_04790_ ), .A2(_04599_ ), .A3(_04562_ ), .ZN(_05196_ ) );
OAI21_X1 _12531_ ( .A(_04899_ ), .B1(_04779_ ), .B2(_04775_ ), .ZN(_05197_ ) );
OAI21_X1 _12532_ ( .A(_04615_ ), .B1(_04768_ ), .B2(_04775_ ), .ZN(_05198_ ) );
OR3_X1 _12533_ ( .A1(_04481_ ), .A2(_03413_ ), .A3(_04487_ ), .ZN(_05199_ ) );
OR2_X1 _12534_ ( .A1(_04493_ ), .A2(_04484_ ), .ZN(_05200_ ) );
OAI21_X1 _12535_ ( .A(_05199_ ), .B1(fanout_net_16 ), .B2(_05200_ ), .ZN(_05201_ ) );
MUX2_X1 _12536_ ( .A(_05126_ ), .B(_05201_ ), .S(_03455_ ), .Z(_05202_ ) );
MUX2_X1 _12537_ ( .A(_05026_ ), .B(_05202_ ), .S(_04518_ ), .Z(_05203_ ) );
OAI211_X1 _12538_ ( .A(_05197_ ), .B(_05198_ ), .C1(_05203_ ), .C2(\u_exu.alu_p2[4] ), .ZN(_05204_ ) );
AOI221_X4 _12539_ ( .A(_05196_ ), .B1(_03112_ ), .B2(_04573_ ), .C1(_05204_ ), .C2(_04717_ ), .ZN(_05205_ ) );
NOR2_X1 _12540_ ( .A1(_03232_ ), .A2(_03234_ ), .ZN(_05206_ ) );
INV_X1 _12541_ ( .A(_03226_ ), .ZN(_05207_ ) );
NOR2_X1 _12542_ ( .A1(_05206_ ), .A2(_05207_ ), .ZN(_05208_ ) );
OR3_X1 _12543_ ( .A1(_05208_ ), .A2(_03222_ ), .A3(_03236_ ), .ZN(_05209_ ) );
OAI21_X1 _12544_ ( .A(_03222_ ), .B1(_05208_ ), .B2(_03236_ ), .ZN(_05210_ ) );
NAND3_X1 _12545_ ( .A1(_05209_ ), .A2(_04478_ ), .A3(_05210_ ), .ZN(_05211_ ) );
OAI211_X1 _12546_ ( .A(_04915_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p2[3] ), .C2(\u_exu.alu_p1[3] ), .ZN(_05212_ ) );
AOI21_X1 _12547_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p2[3] ), .B2(\u_exu.alu_p1[3] ), .ZN(_05213_ ) );
OR2_X1 _12548_ ( .A1(_05212_ ), .A2(_05213_ ), .ZN(_05214_ ) );
NAND4_X1 _12549_ ( .A1(_05205_ ), .A2(_05211_ ), .A3(_04577_ ), .A4(_05214_ ), .ZN(_05215_ ) );
OAI21_X1 _12550_ ( .A(_05215_ ), .B1(\u_exu.alu_p1[3] ), .B2(_04578_ ), .ZN(_05216_ ) );
NOR2_X1 _12551_ ( .A1(_05216_ ), .A2(_04475_ ), .ZN(_00325_ ) );
AND4_X1 _12552_ ( .A1(_03225_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05217_ ) );
OAI211_X1 _12553_ ( .A(_04915_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_ctrl[0] ), .C2(_03088_ ), .ZN(_05218_ ) );
OAI211_X1 _12554_ ( .A(_03083_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(_04498_ ), .C2(_03225_ ), .ZN(_05219_ ) );
AOI21_X1 _12555_ ( .A(_03089_ ), .B1(_05218_ ), .B2(_05219_ ), .ZN(_05220_ ) );
OAI21_X1 _12556_ ( .A(_04478_ ), .B1(_05206_ ), .B2(_05207_ ), .ZN(_05221_ ) );
AOI21_X1 _12557_ ( .A(_05221_ ), .B1(_05206_ ), .B2(_05207_ ), .ZN(_05222_ ) );
OAI21_X1 _12558_ ( .A(_04615_ ), .B1(_04821_ ), .B2(_04828_ ), .ZN(_05223_ ) );
OAI21_X1 _12559_ ( .A(_04899_ ), .B1(_04830_ ), .B2(_04828_ ), .ZN(_05224_ ) );
OR3_X1 _12560_ ( .A1(_03428_ ), .A2(_03429_ ), .A3(_04528_ ), .ZN(_05225_ ) );
OAI211_X1 _12561_ ( .A(_05225_ ), .B(_04498_ ), .C1(\u_exu.alu_p2[1] ), .C2(_03423_ ), .ZN(_05226_ ) );
NAND3_X1 _12562_ ( .A1(_05146_ ), .A2(_05147_ ), .A3(\u_exu.alu_p2[2] ), .ZN(_05227_ ) );
AND3_X1 _12563_ ( .A1(_05226_ ), .A2(_04520_ ), .A3(_05227_ ), .ZN(_05228_ ) );
OAI21_X1 _12564_ ( .A(_04679_ ), .B1(_05051_ ), .B2(_04524_ ), .ZN(_05229_ ) );
OAI211_X1 _12565_ ( .A(_05223_ ), .B(_05224_ ), .C1(_05228_ ), .C2(_05229_ ), .ZN(_05230_ ) );
AOI211_X1 _12566_ ( .A(_05220_ ), .B(_05222_ ), .C1(_04717_ ), .C2(_05230_ ), .ZN(_05231_ ) );
NAND3_X1 _12567_ ( .A1(_04807_ ), .A2(_04524_ ), .A3(_04563_ ), .ZN(_05232_ ) );
AND2_X1 _12568_ ( .A1(_05232_ ), .A2(_04577_ ), .ZN(_05233_ ) );
AOI211_X1 _12569_ ( .A(_04451_ ), .B(_05217_ ), .C1(_05231_ ), .C2(_05233_ ), .ZN(_00326_ ) );
AND4_X1 _12570_ ( .A1(_03351_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05234_ ) );
AOI21_X1 _12571_ ( .A(_04713_ ), .B1(_03344_ ), .B2(_03352_ ), .ZN(_05235_ ) );
OAI21_X1 _12572_ ( .A(_05235_ ), .B1(_03344_ ), .B2(_03352_ ), .ZN(_05236_ ) );
MUX2_X1 _12573_ ( .A(_03361_ ), .B(_04980_ ), .S(_04679_ ), .Z(_05237_ ) );
OR3_X1 _12574_ ( .A1(_05237_ ), .A2(_04982_ ), .A3(_05032_ ), .ZN(_05238_ ) );
OR3_X1 _12575_ ( .A1(_03408_ ), .A2(_03400_ ), .A3(\u_exu.alu_p2[1] ), .ZN(_05239_ ) );
OAI211_X1 _12576_ ( .A(_03405_ ), .B(\u_exu.alu_p2[1] ), .C1(\u_exu.alu_p2[0] ), .C2(_03321_ ), .ZN(_05240_ ) );
NAND3_X1 _12577_ ( .A1(_05239_ ), .A2(_05240_ ), .A3(_04490_ ), .ZN(_05241_ ) );
OR3_X1 _12578_ ( .A1(_04633_ ), .A2(_03392_ ), .A3(_04496_ ), .ZN(_05242_ ) );
NAND3_X1 _12579_ ( .A1(_03403_ ), .A2(_04502_ ), .A3(_03395_ ), .ZN(_05243_ ) );
NAND2_X1 _12580_ ( .A1(_05242_ ), .A2(_05243_ ), .ZN(_05244_ ) );
OAI211_X1 _12581_ ( .A(_05241_ ), .B(_04523_ ), .C1(_05244_ ), .C2(_04498_ ), .ZN(_05245_ ) );
NAND3_X1 _12582_ ( .A1(_04740_ ), .A2(_04743_ ), .A3(\u_exu.alu_p2[3] ), .ZN(_05246_ ) );
AND3_X1 _12583_ ( .A1(_05245_ ), .A2(_05246_ ), .A3(_04679_ ), .ZN(_05247_ ) );
NAND2_X1 _12584_ ( .A1(_05247_ ), .A2(_03378_ ), .ZN(_05248_ ) );
NAND3_X1 _12585_ ( .A1(_04970_ ), .A2(_04501_ ), .A3(_04971_ ), .ZN(_05249_ ) );
OAI211_X1 _12586_ ( .A(_04565_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[28] ), .C2(\u_exu.alu_p2[28] ), .ZN(_05250_ ) );
NAND2_X1 _12587_ ( .A1(\u_exu.alu_p1[28] ), .A2(\u_exu.alu_p2[28] ), .ZN(_05251_ ) );
AOI21_X1 _12588_ ( .A(_05250_ ), .B1(_04962_ ), .B2(_05251_ ), .ZN(_05252_ ) );
AOI211_X1 _12589_ ( .A(_03070_ ), .B(_05252_ ), .C1(_03099_ ), .C2(_04574_ ), .ZN(_05253_ ) );
AND4_X1 _12590_ ( .A1(_05238_ ), .A2(_05248_ ), .A3(_05249_ ), .A4(_05253_ ), .ZN(_05254_ ) );
AOI211_X1 _12591_ ( .A(_04451_ ), .B(_05234_ ), .C1(_05236_ ), .C2(_05254_ ), .ZN(_00327_ ) );
OAI21_X1 _12592_ ( .A(_04615_ ), .B1(_04849_ ), .B2(_04844_ ), .ZN(_05255_ ) );
OAI21_X1 _12593_ ( .A(_04899_ ), .B1(_04839_ ), .B2(_04844_ ), .ZN(_05256_ ) );
NOR3_X1 _12594_ ( .A1(_05077_ ), .A2(_05078_ ), .A3(_04523_ ), .ZN(_05257_ ) );
INV_X1 _12595_ ( .A(_04494_ ), .ZN(_05258_ ) );
AOI21_X1 _12596_ ( .A(\u_exu.alu_p2[1] ), .B1(_05258_ ), .B2(_04700_ ), .ZN(_05259_ ) );
AOI211_X1 _12597_ ( .A(\u_exu.alu_p2[2] ), .B(_05259_ ), .C1(\u_exu.alu_p2[1] ), .C2(_05200_ ), .ZN(_05260_ ) );
AOI21_X1 _12598_ ( .A(_05260_ ), .B1(\u_exu.alu_p2[2] ), .B2(_05169_ ), .ZN(_05261_ ) );
AOI21_X1 _12599_ ( .A(_05257_ ), .B1(_05261_ ), .B2(_04520_ ), .ZN(_05262_ ) );
OAI211_X1 _12600_ ( .A(_05255_ ), .B(_05256_ ), .C1(\u_exu.alu_p2[4] ), .C2(_05262_ ), .ZN(_05263_ ) );
NAND2_X1 _12601_ ( .A1(_05263_ ), .A2(_04717_ ), .ZN(_05264_ ) );
AOI21_X1 _12602_ ( .A(_03229_ ), .B1(_03230_ ), .B2(_03231_ ), .ZN(_05265_ ) );
OR3_X1 _12603_ ( .A1(_03232_ ), .A2(_05265_ ), .A3(_04713_ ), .ZN(_05266_ ) );
OAI211_X1 _12604_ ( .A(_04642_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p2[1] ), .C2(\u_exu.alu_p1[1] ), .ZN(_05267_ ) );
AOI21_X1 _12605_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p2[1] ), .B2(\u_exu.alu_p1[1] ), .ZN(_05268_ ) );
NOR2_X1 _12606_ ( .A1(_05267_ ), .A2(_05268_ ), .ZN(_05269_ ) );
AND4_X1 _12607_ ( .A1(_04600_ ), .A2(_04637_ ), .A3(_04498_ ), .A4(_04701_ ), .ZN(_05270_ ) );
AOI211_X1 _12608_ ( .A(_05269_ ), .B(_05270_ ), .C1(_03086_ ), .C2(_04574_ ), .ZN(_05271_ ) );
AND4_X1 _12609_ ( .A1(_04577_ ), .A2(_05264_ ), .A3(_05266_ ), .A4(_05271_ ), .ZN(_05272_ ) );
NOR4_X1 _12610_ ( .A1(_03379_ ), .A2(\u_exu.alu_p1[1] ), .A3(\u_exu.alu_ctrl[5] ), .A4(\u_exu.alu_ctrl[4] ), .ZN(_05273_ ) );
NOR3_X1 _12611_ ( .A1(_05272_ ), .A2(_01076_ ), .A3(_05273_ ), .ZN(_00328_ ) );
AND3_X1 _12612_ ( .A1(_03467_ ), .A2(_04468_ ), .A3(_03468_ ), .ZN(_00329_ ) );
NAND2_X1 _12613_ ( .A1(_03314_ ), .A2(_03331_ ), .ZN(_05274_ ) );
AOI21_X1 _12614_ ( .A(_03337_ ), .B1(_05274_ ), .B2(_03335_ ), .ZN(_05275_ ) );
NOR3_X1 _12615_ ( .A1(_05275_ ), .A2(_03318_ ), .A3(_03340_ ), .ZN(_05276_ ) );
NOR2_X1 _12616_ ( .A1(_05276_ ), .A2(_04712_ ), .ZN(_05277_ ) );
OAI21_X1 _12617_ ( .A(_03318_ ), .B1(_05275_ ), .B2(_03340_ ), .ZN(_05278_ ) );
AND2_X1 _12618_ ( .A1(_05277_ ), .A2(_05278_ ), .ZN(_05279_ ) );
AND2_X1 _12619_ ( .A1(\u_exu.alu_p1[31] ), .A2(\u_exu.alu_p2[4] ), .ZN(_05280_ ) );
INV_X1 _12620_ ( .A(_05280_ ), .ZN(_05281_ ) );
OAI21_X1 _12621_ ( .A(_05281_ ), .B1(_05030_ ), .B2(\u_exu.alu_p2[4] ), .ZN(_05282_ ) );
NAND2_X1 _12622_ ( .A1(_04778_ ), .A2(_04519_ ), .ZN(_05283_ ) );
AOI21_X1 _12623_ ( .A(_05032_ ), .B1(_05283_ ), .B2(_03366_ ), .ZN(_05284_ ) );
AND2_X1 _12624_ ( .A1(_05282_ ), .A2(_05284_ ), .ZN(_05285_ ) );
OAI211_X1 _12625_ ( .A(_04565_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[27] ), .C2(\u_exu.alu_p2[27] ), .ZN(_05286_ ) );
NAND2_X1 _12626_ ( .A1(\u_exu.alu_p1[27] ), .A2(\u_exu.alu_p2[27] ), .ZN(_05287_ ) );
AOI21_X1 _12627_ ( .A(_05286_ ), .B1(_04962_ ), .B2(_05287_ ), .ZN(_05288_ ) );
AOI21_X1 _12628_ ( .A(_04519_ ), .B1(_04786_ ), .B2(_04787_ ), .ZN(_05289_ ) );
NAND3_X1 _12629_ ( .A1(_04554_ ), .A2(\u_exu.alu_p2[2] ), .A3(_04559_ ), .ZN(_05290_ ) );
NAND3_X1 _12630_ ( .A1(_04536_ ), .A2(_04541_ ), .A3(_03457_ ), .ZN(_05291_ ) );
AOI21_X1 _12631_ ( .A(\u_exu.alu_p2[3] ), .B1(_05290_ ), .B2(_05291_ ), .ZN(_05292_ ) );
OAI21_X1 _12632_ ( .A(_04562_ ), .B1(_05289_ ), .B2(_05292_ ), .ZN(_05293_ ) );
NAND3_X1 _12633_ ( .A1(_05035_ ), .A2(_05036_ ), .A3(_04500_ ), .ZN(_05294_ ) );
NAND2_X1 _12634_ ( .A1(_03126_ ), .A2(_04573_ ), .ZN(_05295_ ) );
NAND3_X1 _12635_ ( .A1(_05293_ ), .A2(_05294_ ), .A3(_05295_ ), .ZN(_05296_ ) );
OR4_X1 _12636_ ( .A1(_05279_ ), .A2(_05285_ ), .A3(_05288_ ), .A4(_05296_ ), .ZN(_05297_ ) );
MUX2_X1 _12637_ ( .A(\u_exu.alu_p1[27] ), .B(_05297_ ), .S(_04578_ ), .Z(_05298_ ) );
AND2_X1 _12638_ ( .A1(_05298_ ), .A2(_04580_ ), .ZN(_00330_ ) );
AND3_X1 _12639_ ( .A1(_05274_ ), .A2(_03337_ ), .A3(_03335_ ), .ZN(_05299_ ) );
NOR3_X1 _12640_ ( .A1(_05299_ ), .A2(_05275_ ), .A3(_04713_ ), .ZN(_05300_ ) );
OAI211_X1 _12641_ ( .A(_04642_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[26] ), .C2(\u_exu.alu_p2[26] ), .ZN(_05301_ ) );
AOI21_X1 _12642_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[26] ), .B2(\u_exu.alu_p2[26] ), .ZN(_05302_ ) );
NOR2_X1 _12643_ ( .A1(_05301_ ), .A2(_05302_ ), .ZN(_05303_ ) );
AND2_X1 _12644_ ( .A1(_03097_ ), .A2(_04573_ ), .ZN(_05304_ ) );
AOI21_X1 _12645_ ( .A(_04489_ ), .B1(_04632_ ), .B2(_04634_ ), .ZN(_05305_ ) );
AOI21_X1 _12646_ ( .A(\u_exu.alu_p2[2] ), .B1(_04624_ ), .B2(_04625_ ), .ZN(_05306_ ) );
OAI21_X1 _12647_ ( .A(_04519_ ), .B1(_05305_ ), .B2(_05306_ ), .ZN(_05307_ ) );
OAI21_X1 _12648_ ( .A(\u_exu.alu_p2[3] ), .B1(_04803_ ), .B2(_04804_ ), .ZN(_05308_ ) );
NAND3_X1 _12649_ ( .A1(_05307_ ), .A2(_05308_ ), .A3(_04562_ ), .ZN(_05309_ ) );
NAND3_X1 _12650_ ( .A1(_05059_ ), .A2(_04500_ ), .A3(_05060_ ), .ZN(_05310_ ) );
MUX2_X1 _12651_ ( .A(_03361_ ), .B(_05057_ ), .S(_03418_ ), .Z(_05311_ ) );
OAI21_X1 _12652_ ( .A(_04998_ ), .B1(_05053_ ), .B2(\u_exu.alu_ctrl[1] ), .ZN(_05312_ ) );
OAI211_X1 _12653_ ( .A(_05309_ ), .B(_05310_ ), .C1(_05311_ ), .C2(_05312_ ), .ZN(_05313_ ) );
OR4_X1 _12654_ ( .A1(_05300_ ), .A2(_05303_ ), .A3(_05304_ ), .A4(_05313_ ), .ZN(_05314_ ) );
MUX2_X1 _12655_ ( .A(\u_exu.alu_p1[26] ), .B(_05314_ ), .S(_04578_ ), .Z(_05315_ ) );
AND2_X1 _12656_ ( .A1(_05315_ ), .A2(_04580_ ), .ZN(_00331_ ) );
NOR2_X1 _12657_ ( .A1(_03324_ ), .A2(\u_exu.alu_p1[24] ), .ZN(_05316_ ) );
NOR3_X1 _12658_ ( .A1(_03313_ ), .A2(_03333_ ), .A3(_05316_ ), .ZN(_05317_ ) );
OR3_X1 _12659_ ( .A1(_05317_ ), .A2(_03333_ ), .A3(_03330_ ), .ZN(_05318_ ) );
OAI21_X1 _12660_ ( .A(_03330_ ), .B1(_05317_ ), .B2(_03333_ ), .ZN(_05319_ ) );
AND3_X1 _12661_ ( .A1(_05318_ ), .A2(_04478_ ), .A3(_05319_ ), .ZN(_05320_ ) );
OAI211_X1 _12662_ ( .A(_04565_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[25] ), .C2(\u_exu.alu_p2[25] ), .ZN(_05321_ ) );
NAND2_X1 _12663_ ( .A1(\u_exu.alu_p1[25] ), .A2(\u_exu.alu_p2[25] ), .ZN(_05322_ ) );
AOI21_X1 _12664_ ( .A(_05321_ ), .B1(_04962_ ), .B2(_05322_ ), .ZN(_05323_ ) );
AND2_X1 _12665_ ( .A1(_04639_ ), .A2(_03100_ ), .ZN(_05324_ ) );
OAI21_X1 _12666_ ( .A(_03418_ ), .B1(_05071_ ), .B2(_04613_ ), .ZN(_05325_ ) );
AOI21_X1 _12667_ ( .A(_03366_ ), .B1(_05325_ ), .B2(_05281_ ), .ZN(_05326_ ) );
NOR4_X1 _12668_ ( .A1(_04838_ ), .A2(\u_exu.alu_ctrl[1] ), .A3(\u_exu.alu_p2[4] ), .A4(\u_exu.alu_p2[3] ), .ZN(_05327_ ) );
OAI21_X1 _12669_ ( .A(_03380_ ), .B1(_05326_ ), .B2(_05327_ ), .ZN(_05328_ ) );
NAND3_X1 _12670_ ( .A1(_05086_ ), .A2(_04500_ ), .A3(_05087_ ), .ZN(_05329_ ) );
AOI21_X1 _12671_ ( .A(_04599_ ), .B1(_04852_ ), .B2(_04853_ ), .ZN(_05330_ ) );
NAND3_X1 _12672_ ( .A1(_04695_ ), .A2(_04696_ ), .A3(\u_exu.alu_p2[2] ), .ZN(_05331_ ) );
NAND3_X1 _12673_ ( .A1(_05001_ ), .A2(_05002_ ), .A3(_04489_ ), .ZN(_05332_ ) );
AOI21_X1 _12674_ ( .A(\u_exu.alu_p2[3] ), .B1(_05331_ ), .B2(_05332_ ), .ZN(_05333_ ) );
OAI21_X1 _12675_ ( .A(_04562_ ), .B1(_05330_ ), .B2(_05333_ ), .ZN(_05334_ ) );
NAND3_X1 _12676_ ( .A1(_05328_ ), .A2(_05329_ ), .A3(_05334_ ), .ZN(_05335_ ) );
OR4_X1 _12677_ ( .A1(_05320_ ), .A2(_05323_ ), .A3(_05324_ ), .A4(_05335_ ), .ZN(_05336_ ) );
MUX2_X1 _12678_ ( .A(\u_exu.alu_p1[25] ), .B(_05336_ ), .S(_04578_ ), .Z(_05337_ ) );
AND2_X1 _12679_ ( .A1(_05337_ ), .A2(_04580_ ), .ZN(_00332_ ) );
AOI21_X1 _12680_ ( .A(_04713_ ), .B1(_03314_ ), .B2(_03326_ ), .ZN(_05338_ ) );
OAI21_X1 _12681_ ( .A(_05338_ ), .B1(_03314_ ), .B2(_03326_ ), .ZN(_05339_ ) );
OAI21_X1 _12682_ ( .A(\u_exu.alu_p2[3] ), .B1(_04871_ ), .B2(_04872_ ), .ZN(_05340_ ) );
NAND2_X1 _12683_ ( .A1(_04739_ ), .A2(\u_exu.alu_p2[2] ), .ZN(_05341_ ) );
OAI211_X1 _12684_ ( .A(_05341_ ), .B(_03454_ ), .C1(\u_exu.alu_p2[2] ), .C2(_05244_ ), .ZN(_05342_ ) );
AND3_X1 _12685_ ( .A1(_05340_ ), .A2(_05342_ ), .A3(_04562_ ), .ZN(_05343_ ) );
INV_X1 _12686_ ( .A(_04500_ ), .ZN(_05344_ ) );
AOI21_X1 _12687_ ( .A(_05344_ ), .B1(_05104_ ), .B2(_05105_ ), .ZN(_05345_ ) );
OR2_X1 _12688_ ( .A1(_05343_ ), .A2(_05345_ ), .ZN(_05346_ ) );
OAI21_X1 _12689_ ( .A(_04998_ ), .B1(_05097_ ), .B2(\u_exu.alu_ctrl[1] ), .ZN(_05347_ ) );
OAI21_X1 _12690_ ( .A(_04679_ ), .B1(_05097_ ), .B2(_04979_ ), .ZN(_05348_ ) );
AOI21_X1 _12691_ ( .A(_05347_ ), .B1(_05281_ ), .B2(_05348_ ), .ZN(_05349_ ) );
AOI211_X1 _12692_ ( .A(_05346_ ), .B(_05349_ ), .C1(_03127_ ), .C2(_04574_ ), .ZN(_05350_ ) );
AOI21_X1 _12693_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[24] ), .B2(\u_exu.alu_p2[24] ), .ZN(_05351_ ) );
OAI211_X1 _12694_ ( .A(_04915_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[24] ), .C2(\u_exu.alu_p2[24] ), .ZN(_05352_ ) );
OAI211_X1 _12695_ ( .A(_05339_ ), .B(_05350_ ), .C1(_05351_ ), .C2(_05352_ ), .ZN(_05353_ ) );
MUX2_X1 _12696_ ( .A(\u_exu.alu_p1[24] ), .B(_05353_ ), .S(_04578_ ), .Z(_05354_ ) );
AND2_X1 _12697_ ( .A1(_05354_ ), .A2(_04580_ ), .ZN(_00333_ ) );
AND4_X1 _12698_ ( .A1(_03265_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05355_ ) );
INV_X1 _12699_ ( .A(_03270_ ), .ZN(_05356_ ) );
NAND2_X1 _12700_ ( .A1(_04714_ ), .A2(_03262_ ), .ZN(_05357_ ) );
AOI21_X1 _12701_ ( .A(_05356_ ), .B1(_05357_ ), .B2(_03307_ ), .ZN(_05358_ ) );
OR3_X1 _12702_ ( .A1(_05358_ ), .A2(_03266_ ), .A3(_03309_ ), .ZN(_05359_ ) );
OAI21_X1 _12703_ ( .A(_03266_ ), .B1(_05358_ ), .B2(_03309_ ), .ZN(_05360_ ) );
NAND3_X1 _12704_ ( .A1(_05359_ ), .A2(_04586_ ), .A3(_05360_ ), .ZN(_05361_ ) );
NOR2_X1 _12705_ ( .A1(_05121_ ), .A2(\u_exu.alu_p2[4] ), .ZN(_05362_ ) );
AOI211_X1 _12706_ ( .A(_03361_ ), .B(_03366_ ), .C1(_04679_ ), .C2(_04520_ ), .ZN(_05363_ ) );
OAI21_X1 _12707_ ( .A(_04717_ ), .B1(_05362_ ), .B2(_05363_ ), .ZN(_05364_ ) );
NAND3_X1 _12708_ ( .A1(_04510_ ), .A2(_04517_ ), .A3(\u_exu.alu_p2[3] ), .ZN(_05365_ ) );
NAND3_X1 _12709_ ( .A1(_04551_ ), .A2(_04560_ ), .A3(_04524_ ), .ZN(_05366_ ) );
NAND3_X1 _12710_ ( .A1(_05365_ ), .A2(_05366_ ), .A3(_04563_ ), .ZN(_05367_ ) );
NAND3_X1 _12711_ ( .A1(_05130_ ), .A2(_04524_ ), .A3(_04501_ ), .ZN(_05368_ ) );
OAI211_X1 _12712_ ( .A(_04565_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[23] ), .C2(\u_exu.alu_p2[23] ), .ZN(_05369_ ) );
NAND2_X1 _12713_ ( .A1(\u_exu.alu_p1[23] ), .A2(\u_exu.alu_p2[23] ), .ZN(_05370_ ) );
AOI21_X1 _12714_ ( .A(_05369_ ), .B1(_04962_ ), .B2(_05370_ ), .ZN(_05371_ ) );
AOI211_X1 _12715_ ( .A(_03070_ ), .B(_05371_ ), .C1(_03123_ ), .C2(_04574_ ), .ZN(_05372_ ) );
AND4_X1 _12716_ ( .A1(_05364_ ), .A2(_05367_ ), .A3(_05368_ ), .A4(_05372_ ), .ZN(_05373_ ) );
AOI211_X1 _12717_ ( .A(_04451_ ), .B(_05355_ ), .C1(_05361_ ), .C2(_05373_ ), .ZN(_00334_ ) );
AND4_X1 _12718_ ( .A1(_03269_ ), .A2(_04583_ ), .A3(_04584_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05374_ ) );
AND3_X1 _12719_ ( .A1(_05357_ ), .A2(_05356_ ), .A3(_03307_ ), .ZN(_05375_ ) );
OR3_X1 _12720_ ( .A1(_05375_ ), .A2(_05358_ ), .A3(_04713_ ), .ZN(_05376_ ) );
OAI21_X1 _12721_ ( .A(_04618_ ), .B1(_05141_ ), .B2(_05142_ ), .ZN(_05377_ ) );
OAI21_X1 _12722_ ( .A(_04609_ ), .B1(_05141_ ), .B2(_05144_ ), .ZN(_05378_ ) );
AND2_X1 _12723_ ( .A1(_05377_ ), .A2(_05378_ ), .ZN(_05379_ ) );
AOI21_X1 _12724_ ( .A(_04571_ ), .B1(_05379_ ), .B2(_04677_ ), .ZN(_05380_ ) );
OAI21_X1 _12725_ ( .A(\u_exu.alu_p2[3] ), .B1(_04603_ ), .B2(_04606_ ), .ZN(_05381_ ) );
NAND3_X1 _12726_ ( .A1(_04631_ ), .A2(_04635_ ), .A3(_04520_ ), .ZN(_05382_ ) );
AND3_X1 _12727_ ( .A1(_05381_ ), .A2(_04563_ ), .A3(_05382_ ), .ZN(_05383_ ) );
AND3_X1 _12728_ ( .A1(_04597_ ), .A2(_04524_ ), .A3(_04501_ ), .ZN(_05384_ ) );
NAND2_X1 _12729_ ( .A1(_03104_ ), .A2(_04639_ ), .ZN(_05385_ ) );
AOI21_X1 _12730_ ( .A(\u_exu.alu_ctrl[0] ), .B1(\u_exu.alu_p1[22] ), .B2(\u_exu.alu_p2[22] ), .ZN(_05386_ ) );
OAI211_X1 _12731_ ( .A(_04642_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1[22] ), .C2(\u_exu.alu_p2[22] ), .ZN(_05387_ ) );
OAI211_X1 _12732_ ( .A(_05385_ ), .B(_03071_ ), .C1(_05386_ ), .C2(_05387_ ), .ZN(_05388_ ) );
NOR4_X1 _12733_ ( .A1(_05380_ ), .A2(_05383_ ), .A3(_05384_ ), .A4(_05388_ ), .ZN(_05389_ ) );
AOI211_X1 _12734_ ( .A(_04451_ ), .B(_05374_ ), .C1(_05376_ ), .C2(_05389_ ), .ZN(_00335_ ) );
BUF_X4 _12735_ ( .A(_00879_ ), .Z(_05390_ ) );
INV_X1 _12736_ ( .A(\fc_addr[31] ), .ZN(_05391_ ) );
NOR3_X1 _12737_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05391_ ), .ZN(_00336_ ) );
BUF_X2 _12738_ ( .A(_01230_ ), .Z(_05392_ ) );
AND3_X1 _12739_ ( .A1(_01226_ ), .A2(_01235_ ), .A3(_01239_ ), .ZN(_05393_ ) );
AND3_X1 _12740_ ( .A1(_01223_ ), .A2(_05392_ ), .A3(_05393_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ) );
CLKBUF_X2 _12741_ ( .A(_00673_ ), .Z(_05394_ ) );
AND4_X1 _12742_ ( .A1(_05394_ ), .A2(_01064_ ), .A3(_01067_ ), .A4(_00968_ ), .ZN(_05395_ ) );
OAI21_X1 _12743_ ( .A(_04468_ ), .B1(_05395_ ), .B2(\u_exu.rlock[15] ), .ZN(_05396_ ) );
NOR2_X1 _12744_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ), .A2(_05396_ ), .ZN(_00337_ ) );
BUF_X2 _12745_ ( .A(_01060_ ), .Z(_05397_ ) );
NAND2_X1 _12746_ ( .A1(_01077_ ), .A2(_00673_ ), .ZN(_05398_ ) );
NOR3_X1 _12747_ ( .A1(_05398_ ), .A2(_00960_ ), .A3(_00942_ ), .ZN(_05399_ ) );
OAI21_X1 _12748_ ( .A(_05397_ ), .B1(_05399_ ), .B2(\u_exu.rlock[14] ), .ZN(_05400_ ) );
INV_X1 _12749_ ( .A(_01226_ ), .ZN(_05401_ ) );
AND3_X1 _12750_ ( .A1(_05401_ ), .A2(_01235_ ), .A3(_01239_ ), .ZN(_05402_ ) );
AND3_X1 _12751_ ( .A1(_01223_ ), .A2(_05392_ ), .A3(_05402_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _12752_ ( .A1(_05400_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_00338_ ) );
AND4_X1 _12753_ ( .A1(_05394_ ), .A2(_01064_ ), .A3(_01067_ ), .A4(_01001_ ), .ZN(_05403_ ) );
OAI21_X1 _12754_ ( .A(_05397_ ), .B1(_05403_ ), .B2(\u_exu.rlock[5] ), .ZN(_05404_ ) );
INV_X1 _12755_ ( .A(_01235_ ), .ZN(_05405_ ) );
AND3_X1 _12756_ ( .A1(_05405_ ), .A2(_01226_ ), .A3(_01239_ ), .ZN(_05406_ ) );
INV_X1 _12757_ ( .A(_05406_ ), .ZN(_05407_ ) );
AOI211_X1 _12758_ ( .A(_05392_ ), .B(_05407_ ), .C1(_01218_ ), .C2(_01220_ ), .ZN(_05408_ ) );
NOR2_X1 _12759_ ( .A1(_05404_ ), .A2(_05408_ ), .ZN(_00339_ ) );
NAND3_X1 _12760_ ( .A1(_05401_ ), .A2(_05405_ ), .A3(_01239_ ), .ZN(_05409_ ) );
NOR3_X1 _12761_ ( .A1(_01222_ ), .A2(_05392_ ), .A3(_05409_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ) );
BUF_X4 _12762_ ( .A(_01060_ ), .Z(_05410_ ) );
AND4_X1 _12763_ ( .A1(_05394_ ), .A2(_01064_ ), .A3(_01041_ ), .A4(_01066_ ), .ZN(_05411_ ) );
OAI21_X1 _12764_ ( .A(_05410_ ), .B1(_05411_ ), .B2(\u_exu.rlock[4] ), .ZN(_05412_ ) );
NOR2_X1 _12765_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ), .A2(_05412_ ), .ZN(_00340_ ) );
AND3_X1 _12766_ ( .A1(_01240_ ), .A2(_01226_ ), .A3(_01235_ ), .ZN(_05413_ ) );
INV_X1 _12767_ ( .A(_05413_ ), .ZN(_05414_ ) );
NOR3_X1 _12768_ ( .A1(_01222_ ), .A2(_05392_ ), .A3(_05414_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ) );
AND4_X1 _12769_ ( .A1(_05394_ ), .A2(_01064_ ), .A3(_01067_ ), .A4(_01013_ ), .ZN(_05415_ ) );
OAI21_X1 _12770_ ( .A(_05410_ ), .B1(_05415_ ), .B2(\u_exu.rlock[3] ), .ZN(_05416_ ) );
NOR2_X1 _12771_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ), .A2(_05416_ ), .ZN(_00341_ ) );
NOR3_X1 _12772_ ( .A1(_05398_ ), .A2(_00946_ ), .A3(_00974_ ), .ZN(_05417_ ) );
OAI21_X1 _12773_ ( .A(_05397_ ), .B1(_05417_ ), .B2(\u_exu.rlock[2] ), .ZN(_05418_ ) );
NOR3_X1 _12774_ ( .A1(_05405_ ), .A2(_01226_ ), .A3(_01239_ ), .ZN(_05419_ ) );
INV_X1 _12775_ ( .A(_05419_ ), .ZN(_05420_ ) );
NOR3_X1 _12776_ ( .A1(_01222_ ), .A2(_05392_ ), .A3(_05420_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _12777_ ( .A1(_05418_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_00342_ ) );
NOR3_X1 _12778_ ( .A1(_05398_ ), .A2(_00946_ ), .A3(_01007_ ), .ZN(_05421_ ) );
OAI21_X1 _12779_ ( .A(_05397_ ), .B1(_05421_ ), .B2(\u_exu.rlock[1] ), .ZN(_05422_ ) );
NOR3_X1 _12780_ ( .A1(_05401_ ), .A2(_01235_ ), .A3(_01239_ ), .ZN(_05423_ ) );
INV_X1 _12781_ ( .A(_05423_ ), .ZN(_05424_ ) );
AOI211_X1 _12782_ ( .A(_05392_ ), .B(_05424_ ), .C1(_01218_ ), .C2(_01220_ ), .ZN(_05425_ ) );
NOR2_X1 _12783_ ( .A1(_05422_ ), .A2(_05425_ ), .ZN(_00343_ ) );
NOR3_X1 _12784_ ( .A1(_01226_ ), .A2(_01235_ ), .A3(_01239_ ), .ZN(_05426_ ) );
INV_X1 _12785_ ( .A(_05426_ ), .ZN(_05427_ ) );
NOR3_X1 _12786_ ( .A1(_01222_ ), .A2(_05392_ ), .A3(_05427_ ), .ZN(_05428_ ) );
AND4_X1 _12787_ ( .A1(_05394_ ), .A2(_01064_ ), .A3(_01067_ ), .A4(_00985_ ), .ZN(_05429_ ) );
OAI21_X1 _12788_ ( .A(_05410_ ), .B1(_05429_ ), .B2(\u_exu.rlock[0] ), .ZN(_05430_ ) );
NOR2_X1 _12789_ ( .A1(_05428_ ), .A2(_05430_ ), .ZN(_00344_ ) );
NOR3_X1 _12790_ ( .A1(_01222_ ), .A2(_01231_ ), .A3(_05407_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ) );
AND4_X1 _12791_ ( .A1(_05394_ ), .A2(_01064_ ), .A3(_01067_ ), .A4(_01017_ ), .ZN(_05431_ ) );
OAI21_X1 _12792_ ( .A(_05410_ ), .B1(_05431_ ), .B2(\u_exu.rlock[13] ), .ZN(_05432_ ) );
NOR2_X1 _12793_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .A2(_05432_ ), .ZN(_00345_ ) );
NOR3_X1 _12794_ ( .A1(_01222_ ), .A2(_01231_ ), .A3(_05409_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ) );
AND4_X1 _12795_ ( .A1(_05394_ ), .A2(_01063_ ), .A3(_01067_ ), .A4(_00993_ ), .ZN(_05433_ ) );
OAI21_X1 _12796_ ( .A(_05410_ ), .B1(_05433_ ), .B2(\u_exu.rlock[12] ), .ZN(_05434_ ) );
NOR2_X1 _12797_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ), .A2(_05434_ ), .ZN(_00346_ ) );
NOR3_X1 _12798_ ( .A1(_01222_ ), .A2(_01231_ ), .A3(_05414_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ) );
AND4_X1 _12799_ ( .A1(_05394_ ), .A2(_01063_ ), .A3(_01066_ ), .A4(_00961_ ), .ZN(_05435_ ) );
OAI21_X1 _12800_ ( .A(_05410_ ), .B1(_05435_ ), .B2(\u_exu.rlock[11] ), .ZN(_05436_ ) );
NOR2_X1 _12801_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ), .A2(_05436_ ), .ZN(_00347_ ) );
NOR3_X1 _12802_ ( .A1(_05398_ ), .A2(_00960_ ), .A3(_00974_ ), .ZN(_05437_ ) );
OAI21_X1 _12803_ ( .A(_05397_ ), .B1(_05437_ ), .B2(\u_exu.rlock[10] ), .ZN(_05438_ ) );
NOR3_X1 _12804_ ( .A1(_01222_ ), .A2(_01231_ ), .A3(_05420_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _12805_ ( .A1(_05438_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ), .ZN(_00348_ ) );
NOR3_X1 _12806_ ( .A1(_01222_ ), .A2(_01231_ ), .A3(_05424_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ) );
AND4_X1 _12807_ ( .A1(_05394_ ), .A2(_01063_ ), .A3(_01029_ ), .A4(_01066_ ), .ZN(_05439_ ) );
OAI21_X1 _12808_ ( .A(_05410_ ), .B1(_05439_ ), .B2(\u_exu.rlock[9] ), .ZN(_05440_ ) );
NOR2_X1 _12809_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ), .A2(_05440_ ), .ZN(_00349_ ) );
AND4_X1 _12810_ ( .A1(_05394_ ), .A2(_01064_ ), .A3(_01037_ ), .A4(_01067_ ), .ZN(_05441_ ) );
OAI21_X1 _12811_ ( .A(_05397_ ), .B1(_05441_ ), .B2(\u_exu.rlock[8] ), .ZN(_05442_ ) );
AOI211_X1 _12812_ ( .A(_01231_ ), .B(_05427_ ), .C1(_01218_ ), .C2(_01220_ ), .ZN(_05443_ ) );
NOR2_X1 _12813_ ( .A1(_05442_ ), .A2(_05443_ ), .ZN(_00350_ ) );
AND3_X1 _12814_ ( .A1(_01223_ ), .A2(_01231_ ), .A3(_05393_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_Y_$_AND__B_Y ) );
AND4_X1 _12815_ ( .A1(_00673_ ), .A2(_01063_ ), .A3(_01034_ ), .A4(_01066_ ), .ZN(_05444_ ) );
OAI21_X1 _12816_ ( .A(_05410_ ), .B1(_05444_ ), .B2(\u_exu.rlock[7] ), .ZN(_05445_ ) );
NOR2_X1 _12817_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_Y_$_AND__B_Y ), .A2(_05445_ ), .ZN(_00351_ ) );
AND3_X1 _12818_ ( .A1(_01223_ ), .A2(_01231_ ), .A3(_05402_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
AND4_X1 _12819_ ( .A1(_00673_ ), .A2(_01063_ ), .A3(_01066_ ), .A4(_00947_ ), .ZN(_05446_ ) );
OAI21_X1 _12820_ ( .A(_05410_ ), .B1(_05446_ ), .B2(\u_exu.rlock[6] ), .ZN(_05447_ ) );
NOR2_X1 _12821_ ( .A1(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .A2(_05447_ ), .ZN(_00352_ ) );
INV_X1 _12822_ ( .A(\fc_addr[30] ), .ZN(_05448_ ) );
NOR3_X1 _12823_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05448_ ), .ZN(_00353_ ) );
INV_X1 _12824_ ( .A(\fc_addr[21] ), .ZN(_05449_ ) );
NOR3_X1 _12825_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05449_ ), .ZN(_00354_ ) );
INV_X1 _12826_ ( .A(\fc_addr[20] ), .ZN(_05450_ ) );
NOR3_X1 _12827_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05450_ ), .ZN(_00355_ ) );
INV_X1 _12828_ ( .A(\fc_addr[19] ), .ZN(_05451_ ) );
NOR3_X1 _12829_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05451_ ), .ZN(_00356_ ) );
INV_X1 _12830_ ( .A(\fc_addr[18] ), .ZN(_05452_ ) );
NOR3_X1 _12831_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05452_ ), .ZN(_00357_ ) );
INV_X1 _12832_ ( .A(\fc_addr[17] ), .ZN(_05453_ ) );
NOR3_X1 _12833_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05453_ ), .ZN(_00358_ ) );
INV_X1 _12834_ ( .A(\fc_addr[16] ), .ZN(_05454_ ) );
NOR3_X1 _12835_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05454_ ), .ZN(_00359_ ) );
INV_X1 _12836_ ( .A(\fc_addr[15] ), .ZN(_05455_ ) );
NOR3_X1 _12837_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05455_ ), .ZN(_00360_ ) );
INV_X1 _12838_ ( .A(\fc_addr[14] ), .ZN(_05456_ ) );
NOR3_X1 _12839_ ( .A1(_05390_ ), .A2(fanout_net_2 ), .A3(_05456_ ), .ZN(_00361_ ) );
BUF_X4 _12840_ ( .A(_00879_ ), .Z(_05457_ ) );
INV_X1 _12841_ ( .A(\fc_addr[13] ), .ZN(_05458_ ) );
NOR3_X1 _12842_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05458_ ), .ZN(_00362_ ) );
INV_X1 _12843_ ( .A(\fc_addr[12] ), .ZN(_05459_ ) );
NOR3_X1 _12844_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05459_ ), .ZN(_00363_ ) );
INV_X1 _12845_ ( .A(\fc_addr[29] ), .ZN(_05460_ ) );
NOR3_X1 _12846_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05460_ ), .ZN(_00364_ ) );
INV_X1 _12847_ ( .A(\fc_addr[11] ), .ZN(_05461_ ) );
NOR3_X1 _12848_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05461_ ), .ZN(_00365_ ) );
INV_X1 _12849_ ( .A(\fc_addr[10] ), .ZN(_05462_ ) );
NOR3_X1 _12850_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05462_ ), .ZN(_00366_ ) );
INV_X1 _12851_ ( .A(\fc_addr[9] ), .ZN(_05463_ ) );
NOR3_X1 _12852_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05463_ ), .ZN(_00367_ ) );
INV_X1 _12853_ ( .A(\fc_addr[8] ), .ZN(_05464_ ) );
NOR3_X1 _12854_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05464_ ), .ZN(_00368_ ) );
INV_X1 _12855_ ( .A(\fc_addr[7] ), .ZN(_05465_ ) );
NOR3_X1 _12856_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05465_ ), .ZN(_00369_ ) );
INV_X1 _12857_ ( .A(\fc_addr[6] ), .ZN(_05466_ ) );
NOR3_X1 _12858_ ( .A1(_05457_ ), .A2(fanout_net_2 ), .A3(_05466_ ), .ZN(_00370_ ) );
INV_X1 _12859_ ( .A(\fc_addr[5] ), .ZN(_05467_ ) );
NOR3_X1 _12860_ ( .A1(_05457_ ), .A2(fanout_net_3 ), .A3(_05467_ ), .ZN(_00371_ ) );
INV_X1 _12861_ ( .A(fanout_net_10 ), .ZN(_05468_ ) );
BUF_X4 _12862_ ( .A(_05468_ ), .Z(_05469_ ) );
NOR3_X1 _12863_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05469_ ), .ZN(_00372_ ) );
INV_X1 _12864_ ( .A(\fc_addr[28] ), .ZN(_05470_ ) );
NOR3_X1 _12865_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05470_ ), .ZN(_00373_ ) );
INV_X1 _12866_ ( .A(\fc_addr[27] ), .ZN(_05471_ ) );
NOR3_X1 _12867_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05471_ ), .ZN(_00374_ ) );
INV_X1 _12868_ ( .A(\fc_addr[26] ), .ZN(_05472_ ) );
NOR3_X1 _12869_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05472_ ), .ZN(_00375_ ) );
INV_X1 _12870_ ( .A(\fc_addr[25] ), .ZN(_05473_ ) );
NOR3_X1 _12871_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05473_ ), .ZN(_00376_ ) );
INV_X1 _12872_ ( .A(\fc_addr[24] ), .ZN(_05474_ ) );
NOR3_X1 _12873_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05474_ ), .ZN(_00377_ ) );
INV_X1 _12874_ ( .A(\fc_addr[23] ), .ZN(_05475_ ) );
NOR3_X1 _12875_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05475_ ), .ZN(_00378_ ) );
INV_X1 _12876_ ( .A(\fc_addr[22] ), .ZN(_05476_ ) );
NOR3_X1 _12877_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05476_ ), .ZN(_00379_ ) );
INV_X2 _12878_ ( .A(_00863_ ), .ZN(_05477_ ) );
BUF_X4 _12879_ ( .A(_05477_ ), .Z(_05478_ ) );
INV_X1 _12880_ ( .A(fanout_net_6 ), .ZN(_05479_ ) );
BUF_X2 _12881_ ( .A(_05479_ ), .Z(_05480_ ) );
CLKBUF_X2 _12882_ ( .A(_05480_ ), .Z(_05481_ ) );
OR2_X1 _12883_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[1][31] ), .ZN(_05482_ ) );
INV_X1 _12884_ ( .A(fanout_net_8 ), .ZN(_05483_ ) );
BUF_X4 _12885_ ( .A(_05483_ ), .Z(_05484_ ) );
BUF_X4 _12886_ ( .A(_05484_ ), .Z(_05485_ ) );
OR2_X1 _12887_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[0][31] ), .ZN(_05486_ ) );
NAND3_X1 _12888_ ( .A1(_05482_ ), .A2(_05485_ ), .A3(_05486_ ), .ZN(_05487_ ) );
CLKBUF_X2 _12889_ ( .A(_05480_ ), .Z(_05488_ ) );
AND3_X1 _12890_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][31] ), .ZN(_05489_ ) );
AND2_X1 _12891_ ( .A1(fanout_net_8 ), .A2(fanout_net_6 ), .ZN(_05490_ ) );
BUF_X4 _12892_ ( .A(_05490_ ), .Z(_05491_ ) );
BUF_X4 _12893_ ( .A(_05491_ ), .Z(_05492_ ) );
AOI211_X1 _12894_ ( .A(fanout_net_10 ), .B(_05489_ ), .C1(\u_icache.cblocks[3][31] ), .C2(_05492_ ), .ZN(_05493_ ) );
BUF_X4 _12895_ ( .A(_05484_ ), .Z(_05494_ ) );
CLKBUF_X2 _12896_ ( .A(_05480_ ), .Z(_05495_ ) );
CLKBUF_X2 _12897_ ( .A(_05495_ ), .Z(_05496_ ) );
AND2_X1 _12898_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][31] ), .ZN(_05497_ ) );
AND2_X1 _12899_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[5][31] ), .ZN(_05498_ ) );
OAI21_X1 _12900_ ( .A(_05494_ ), .B1(_05497_ ), .B2(_05498_ ), .ZN(_05499_ ) );
CLKBUF_X2 _12901_ ( .A(_05480_ ), .Z(_05500_ ) );
AND3_X1 _12902_ ( .A1(_05500_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][31] ), .ZN(_05501_ ) );
BUF_X4 _12903_ ( .A(_05491_ ), .Z(_05502_ ) );
AOI211_X1 _12904_ ( .A(_05469_ ), .B(_05501_ ), .C1(\u_icache.cblocks[7][31] ), .C2(_05502_ ), .ZN(_05503_ ) );
AOI221_X4 _12905_ ( .A(_05478_ ), .B1(_05487_ ), .B2(_05493_ ), .C1(_05499_ ), .C2(_05503_ ), .ZN(_00380_ ) );
OR2_X1 _12906_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[1][30] ), .ZN(_05504_ ) );
OR2_X1 _12907_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[0][30] ), .ZN(_05505_ ) );
NAND3_X1 _12908_ ( .A1(_05504_ ), .A2(_05485_ ), .A3(_05505_ ), .ZN(_05506_ ) );
AND3_X1 _12909_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][30] ), .ZN(_05507_ ) );
AOI211_X1 _12910_ ( .A(fanout_net_10 ), .B(_05507_ ), .C1(\u_icache.cblocks[3][30] ), .C2(_05492_ ), .ZN(_05508_ ) );
CLKBUF_X2 _12911_ ( .A(_05495_ ), .Z(_05509_ ) );
OR2_X1 _12912_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[5][30] ), .ZN(_05510_ ) );
BUF_X4 _12913_ ( .A(_05484_ ), .Z(_05511_ ) );
OR2_X1 _12914_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[4][30] ), .ZN(_05512_ ) );
NAND3_X1 _12915_ ( .A1(_05510_ ), .A2(_05511_ ), .A3(_05512_ ), .ZN(_05513_ ) );
BUF_X4 _12916_ ( .A(_05468_ ), .Z(_05514_ ) );
AND3_X1 _12917_ ( .A1(_05500_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][30] ), .ZN(_05515_ ) );
AOI211_X1 _12918_ ( .A(_05514_ ), .B(_05515_ ), .C1(\u_icache.cblocks[7][30] ), .C2(_05502_ ), .ZN(_05516_ ) );
AOI221_X4 _12919_ ( .A(_05478_ ), .B1(_05506_ ), .B2(_05508_ ), .C1(_05513_ ), .C2(_05516_ ), .ZN(_00381_ ) );
CLKBUF_X2 _12920_ ( .A(_05480_ ), .Z(_05517_ ) );
OR2_X1 _12921_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][21] ), .ZN(_05518_ ) );
OR2_X1 _12922_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[0][21] ), .ZN(_05519_ ) );
NAND3_X1 _12923_ ( .A1(_05518_ ), .A2(_05485_ ), .A3(_05519_ ), .ZN(_05520_ ) );
AND3_X1 _12924_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][21] ), .ZN(_05521_ ) );
AOI211_X1 _12925_ ( .A(fanout_net_10 ), .B(_05521_ ), .C1(\u_icache.cblocks[3][21] ), .C2(_05492_ ), .ZN(_05522_ ) );
AND2_X1 _12926_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][21] ), .ZN(_05523_ ) );
AND2_X1 _12927_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[5][21] ), .ZN(_05524_ ) );
OAI21_X1 _12928_ ( .A(_05494_ ), .B1(_05523_ ), .B2(_05524_ ), .ZN(_05525_ ) );
AND3_X1 _12929_ ( .A1(_05500_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][21] ), .ZN(_05526_ ) );
AOI211_X1 _12930_ ( .A(_05514_ ), .B(_05526_ ), .C1(\u_icache.cblocks[7][21] ), .C2(_05502_ ), .ZN(_05527_ ) );
AOI221_X4 _12931_ ( .A(_05478_ ), .B1(_05520_ ), .B2(_05522_ ), .C1(_05525_ ), .C2(_05527_ ), .ZN(_00382_ ) );
BUF_X4 _12932_ ( .A(_05483_ ), .Z(_05528_ ) );
CLKBUF_X2 _12933_ ( .A(_05480_ ), .Z(_05529_ ) );
AND2_X1 _12934_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[0][20] ), .ZN(_05530_ ) );
AND2_X1 _12935_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][20] ), .ZN(_05531_ ) );
OAI21_X1 _12936_ ( .A(_05528_ ), .B1(_05530_ ), .B2(_05531_ ), .ZN(_05532_ ) );
AND3_X1 _12937_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][20] ), .ZN(_05533_ ) );
AOI211_X1 _12938_ ( .A(fanout_net_10 ), .B(_05533_ ), .C1(\u_icache.cblocks[3][20] ), .C2(_05492_ ), .ZN(_05534_ ) );
OR2_X1 _12939_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[5][20] ), .ZN(_05535_ ) );
OR2_X1 _12940_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[4][20] ), .ZN(_05536_ ) );
NAND3_X1 _12941_ ( .A1(_05535_ ), .A2(_05511_ ), .A3(_05536_ ), .ZN(_05537_ ) );
AND3_X1 _12942_ ( .A1(_05500_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][20] ), .ZN(_05538_ ) );
AOI211_X1 _12943_ ( .A(_05514_ ), .B(_05538_ ), .C1(\u_icache.cblocks[7][20] ), .C2(_05502_ ), .ZN(_05539_ ) );
AOI221_X4 _12944_ ( .A(_05478_ ), .B1(_05532_ ), .B2(_05534_ ), .C1(_05537_ ), .C2(_05539_ ), .ZN(_00383_ ) );
OR2_X1 _12945_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][19] ), .ZN(_05540_ ) );
OR2_X1 _12946_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[0][19] ), .ZN(_05541_ ) );
NAND3_X1 _12947_ ( .A1(_05540_ ), .A2(_05485_ ), .A3(_05541_ ), .ZN(_05542_ ) );
AND3_X1 _12948_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][19] ), .ZN(_05543_ ) );
AOI211_X1 _12949_ ( .A(fanout_net_10 ), .B(_05543_ ), .C1(\u_icache.cblocks[3][19] ), .C2(_05492_ ), .ZN(_05544_ ) );
BUF_X4 _12950_ ( .A(_05484_ ), .Z(_05545_ ) );
AND2_X1 _12951_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][19] ), .ZN(_05546_ ) );
AND2_X1 _12952_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[5][19] ), .ZN(_05547_ ) );
OAI21_X1 _12953_ ( .A(_05545_ ), .B1(_05546_ ), .B2(_05547_ ), .ZN(_05548_ ) );
AND3_X1 _12954_ ( .A1(_05500_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][19] ), .ZN(_05549_ ) );
AOI211_X1 _12955_ ( .A(_05514_ ), .B(_05549_ ), .C1(\u_icache.cblocks[7][19] ), .C2(_05502_ ), .ZN(_05550_ ) );
AOI221_X4 _12956_ ( .A(_05478_ ), .B1(_05542_ ), .B2(_05544_ ), .C1(_05548_ ), .C2(_05550_ ), .ZN(_00384_ ) );
AND2_X1 _12957_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[0][18] ), .ZN(_05551_ ) );
AND2_X1 _12958_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][18] ), .ZN(_05552_ ) );
OAI21_X1 _12959_ ( .A(_05528_ ), .B1(_05551_ ), .B2(_05552_ ), .ZN(_05553_ ) );
AND3_X1 _12960_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][18] ), .ZN(_05554_ ) );
AOI211_X1 _12961_ ( .A(fanout_net_10 ), .B(_05554_ ), .C1(\u_icache.cblocks[3][18] ), .C2(_05492_ ), .ZN(_05555_ ) );
OR2_X1 _12962_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[5][18] ), .ZN(_05556_ ) );
OR2_X1 _12963_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[4][18] ), .ZN(_05557_ ) );
NAND3_X1 _12964_ ( .A1(_05556_ ), .A2(_05511_ ), .A3(_05557_ ), .ZN(_05558_ ) );
CLKBUF_X2 _12965_ ( .A(_05480_ ), .Z(_05559_ ) );
AND3_X1 _12966_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][18] ), .ZN(_05560_ ) );
AOI211_X1 _12967_ ( .A(_05514_ ), .B(_05560_ ), .C1(\u_icache.cblocks[7][18] ), .C2(_05502_ ), .ZN(_05561_ ) );
AOI221_X4 _12968_ ( .A(_05478_ ), .B1(_05553_ ), .B2(_05555_ ), .C1(_05558_ ), .C2(_05561_ ), .ZN(_00385_ ) );
BUF_X4 _12969_ ( .A(_05477_ ), .Z(_05562_ ) );
AND2_X1 _12970_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[0][17] ), .ZN(_05563_ ) );
AND2_X1 _12971_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][17] ), .ZN(_05564_ ) );
OAI21_X1 _12972_ ( .A(_05528_ ), .B1(_05563_ ), .B2(_05564_ ), .ZN(_05565_ ) );
AND3_X1 _12973_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][17] ), .ZN(_05566_ ) );
AOI211_X1 _12974_ ( .A(fanout_net_10 ), .B(_05566_ ), .C1(\u_icache.cblocks[3][17] ), .C2(_05492_ ), .ZN(_05567_ ) );
OR2_X1 _12975_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[5][17] ), .ZN(_05568_ ) );
OR2_X1 _12976_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[4][17] ), .ZN(_05569_ ) );
NAND3_X1 _12977_ ( .A1(_05568_ ), .A2(_05511_ ), .A3(_05569_ ), .ZN(_05570_ ) );
AND3_X1 _12978_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][17] ), .ZN(_05571_ ) );
AOI211_X1 _12979_ ( .A(_05514_ ), .B(_05571_ ), .C1(\u_icache.cblocks[7][17] ), .C2(_05502_ ), .ZN(_05572_ ) );
AOI221_X4 _12980_ ( .A(_05562_ ), .B1(_05565_ ), .B2(_05567_ ), .C1(_05570_ ), .C2(_05572_ ), .ZN(_00386_ ) );
OR2_X1 _12981_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][16] ), .ZN(_05573_ ) );
OR2_X1 _12982_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[0][16] ), .ZN(_05574_ ) );
NAND3_X1 _12983_ ( .A1(_05573_ ), .A2(_05485_ ), .A3(_05574_ ), .ZN(_05575_ ) );
AND3_X1 _12984_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][16] ), .ZN(_05576_ ) );
BUF_X4 _12985_ ( .A(_05491_ ), .Z(_05577_ ) );
AOI211_X1 _12986_ ( .A(fanout_net_10 ), .B(_05576_ ), .C1(\u_icache.cblocks[3][16] ), .C2(_05577_ ), .ZN(_05578_ ) );
AND2_X1 _12987_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][16] ), .ZN(_05579_ ) );
AND2_X1 _12988_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[5][16] ), .ZN(_05580_ ) );
OAI21_X1 _12989_ ( .A(_05545_ ), .B1(_05579_ ), .B2(_05580_ ), .ZN(_05581_ ) );
AND3_X1 _12990_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][16] ), .ZN(_05582_ ) );
AOI211_X1 _12991_ ( .A(_05514_ ), .B(_05582_ ), .C1(\u_icache.cblocks[7][16] ), .C2(_05502_ ), .ZN(_05583_ ) );
AOI221_X4 _12992_ ( .A(_05562_ ), .B1(_05575_ ), .B2(_05578_ ), .C1(_05581_ ), .C2(_05583_ ), .ZN(_00387_ ) );
AND2_X1 _12993_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[0][15] ), .ZN(_05584_ ) );
AND2_X1 _12994_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][15] ), .ZN(_05585_ ) );
OAI21_X1 _12995_ ( .A(_05528_ ), .B1(_05584_ ), .B2(_05585_ ), .ZN(_05586_ ) );
AND3_X1 _12996_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][15] ), .ZN(_05587_ ) );
AOI211_X1 _12997_ ( .A(fanout_net_10 ), .B(_05587_ ), .C1(\u_icache.cblocks[3][15] ), .C2(_05577_ ), .ZN(_05588_ ) );
AND2_X1 _12998_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][15] ), .ZN(_05589_ ) );
AND2_X1 _12999_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[5][15] ), .ZN(_05590_ ) );
OAI21_X1 _13000_ ( .A(_05545_ ), .B1(_05589_ ), .B2(_05590_ ), .ZN(_05591_ ) );
AND3_X1 _13001_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][15] ), .ZN(_05592_ ) );
AOI211_X1 _13002_ ( .A(_05514_ ), .B(_05592_ ), .C1(\u_icache.cblocks[7][15] ), .C2(_05502_ ), .ZN(_05593_ ) );
AOI221_X4 _13003_ ( .A(_05562_ ), .B1(_05586_ ), .B2(_05588_ ), .C1(_05591_ ), .C2(_05593_ ), .ZN(_00388_ ) );
OR2_X1 _13004_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][14] ), .ZN(_05594_ ) );
OR2_X1 _13005_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[0][14] ), .ZN(_05595_ ) );
NAND3_X1 _13006_ ( .A1(_05594_ ), .A2(_05485_ ), .A3(_05595_ ), .ZN(_05596_ ) );
AND3_X1 _13007_ ( .A1(_05488_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][14] ), .ZN(_05597_ ) );
AOI211_X1 _13008_ ( .A(fanout_net_10 ), .B(_05597_ ), .C1(\u_icache.cblocks[3][14] ), .C2(_05577_ ), .ZN(_05598_ ) );
CLKBUF_X2 _13009_ ( .A(_05495_ ), .Z(_05599_ ) );
OR2_X1 _13010_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][14] ), .ZN(_05600_ ) );
OR2_X1 _13011_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[4][14] ), .ZN(_05601_ ) );
NAND3_X1 _13012_ ( .A1(_05600_ ), .A2(_05511_ ), .A3(_05601_ ), .ZN(_05602_ ) );
AND3_X1 _13013_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][14] ), .ZN(_05603_ ) );
BUF_X4 _13014_ ( .A(_05491_ ), .Z(_05604_ ) );
AOI211_X1 _13015_ ( .A(_05514_ ), .B(_05603_ ), .C1(\u_icache.cblocks[7][14] ), .C2(_05604_ ), .ZN(_05605_ ) );
AOI221_X4 _13016_ ( .A(_05562_ ), .B1(_05596_ ), .B2(_05598_ ), .C1(_05602_ ), .C2(_05605_ ), .ZN(_00389_ ) );
AND2_X1 _13017_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[0][13] ), .ZN(_05606_ ) );
AND2_X1 _13018_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][13] ), .ZN(_05607_ ) );
OAI21_X1 _13019_ ( .A(_05528_ ), .B1(_05606_ ), .B2(_05607_ ), .ZN(_05608_ ) );
CLKBUF_X2 _13020_ ( .A(_05479_ ), .Z(_05609_ ) );
AND3_X1 _13021_ ( .A1(_05609_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][13] ), .ZN(_05610_ ) );
AOI211_X1 _13022_ ( .A(fanout_net_10 ), .B(_05610_ ), .C1(\u_icache.cblocks[3][13] ), .C2(_05577_ ), .ZN(_05611_ ) );
AND2_X1 _13023_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][13] ), .ZN(_05612_ ) );
AND2_X1 _13024_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[5][13] ), .ZN(_05613_ ) );
OAI21_X1 _13025_ ( .A(_05545_ ), .B1(_05612_ ), .B2(_05613_ ), .ZN(_05614_ ) );
AND3_X1 _13026_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][13] ), .ZN(_05615_ ) );
AOI211_X1 _13027_ ( .A(_05514_ ), .B(_05615_ ), .C1(\u_icache.cblocks[7][13] ), .C2(_05604_ ), .ZN(_05616_ ) );
AOI221_X4 _13028_ ( .A(_05562_ ), .B1(_05608_ ), .B2(_05611_ ), .C1(_05614_ ), .C2(_05616_ ), .ZN(_00390_ ) );
AND2_X1 _13029_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[0][12] ), .ZN(_05617_ ) );
AND2_X1 _13030_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][12] ), .ZN(_05618_ ) );
OAI21_X1 _13031_ ( .A(_05528_ ), .B1(_05617_ ), .B2(_05618_ ), .ZN(_05619_ ) );
AND3_X1 _13032_ ( .A1(_05609_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][12] ), .ZN(_05620_ ) );
AOI211_X1 _13033_ ( .A(fanout_net_10 ), .B(_05620_ ), .C1(\u_icache.cblocks[3][12] ), .C2(_05577_ ), .ZN(_05621_ ) );
OR2_X1 _13034_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][12] ), .ZN(_05622_ ) );
OR2_X1 _13035_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[4][12] ), .ZN(_05623_ ) );
NAND3_X1 _13036_ ( .A1(_05622_ ), .A2(_05511_ ), .A3(_05623_ ), .ZN(_05624_ ) );
BUF_X4 _13037_ ( .A(_05468_ ), .Z(_05625_ ) );
AND3_X1 _13038_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][12] ), .ZN(_05626_ ) );
AOI211_X1 _13039_ ( .A(_05625_ ), .B(_05626_ ), .C1(\u_icache.cblocks[7][12] ), .C2(_05604_ ), .ZN(_05627_ ) );
AOI221_X4 _13040_ ( .A(_05562_ ), .B1(_05619_ ), .B2(_05621_ ), .C1(_05624_ ), .C2(_05627_ ), .ZN(_00391_ ) );
AND2_X1 _13041_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[0][29] ), .ZN(_05628_ ) );
AND2_X1 _13042_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][29] ), .ZN(_05629_ ) );
OAI21_X1 _13043_ ( .A(_05528_ ), .B1(_05628_ ), .B2(_05629_ ), .ZN(_05630_ ) );
AND3_X1 _13044_ ( .A1(_05609_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][29] ), .ZN(_05631_ ) );
AOI211_X1 _13045_ ( .A(fanout_net_10 ), .B(_05631_ ), .C1(\u_icache.cblocks[3][29] ), .C2(_05577_ ), .ZN(_05632_ ) );
AND2_X1 _13046_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][29] ), .ZN(_05633_ ) );
AND2_X1 _13047_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[5][29] ), .ZN(_05634_ ) );
OAI21_X1 _13048_ ( .A(_05545_ ), .B1(_05633_ ), .B2(_05634_ ), .ZN(_05635_ ) );
AND3_X1 _13049_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][29] ), .ZN(_05636_ ) );
AOI211_X1 _13050_ ( .A(_05625_ ), .B(_05636_ ), .C1(\u_icache.cblocks[7][29] ), .C2(_05604_ ), .ZN(_05637_ ) );
AOI221_X4 _13051_ ( .A(_05562_ ), .B1(_05630_ ), .B2(_05632_ ), .C1(_05635_ ), .C2(_05637_ ), .ZN(_00392_ ) );
AND2_X1 _13052_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][11] ), .ZN(_05638_ ) );
AND2_X1 _13053_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[1][11] ), .ZN(_05639_ ) );
OAI21_X1 _13054_ ( .A(_05528_ ), .B1(_05638_ ), .B2(_05639_ ), .ZN(_05640_ ) );
AND3_X1 _13055_ ( .A1(_05609_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[2][11] ), .ZN(_05641_ ) );
AOI211_X1 _13056_ ( .A(fanout_net_10 ), .B(_05641_ ), .C1(\u_icache.cblocks[3][11] ), .C2(_05577_ ), .ZN(_05642_ ) );
OR2_X1 _13057_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][11] ), .ZN(_05643_ ) );
OR2_X1 _13058_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[4][11] ), .ZN(_05644_ ) );
NAND3_X1 _13059_ ( .A1(_05643_ ), .A2(_05511_ ), .A3(_05644_ ), .ZN(_05645_ ) );
AND3_X1 _13060_ ( .A1(_05559_ ), .A2(fanout_net_8 ), .A3(\u_icache.cblocks[6][11] ), .ZN(_05646_ ) );
AOI211_X1 _13061_ ( .A(_05625_ ), .B(_05646_ ), .C1(\u_icache.cblocks[7][11] ), .C2(_05604_ ), .ZN(_05647_ ) );
AOI221_X4 _13062_ ( .A(_05562_ ), .B1(_05640_ ), .B2(_05642_ ), .C1(_05645_ ), .C2(_05647_ ), .ZN(_00393_ ) );
OR2_X1 _13063_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][10] ), .ZN(_05648_ ) );
OR2_X1 _13064_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][10] ), .ZN(_05649_ ) );
NAND3_X1 _13065_ ( .A1(_05648_ ), .A2(_05485_ ), .A3(_05649_ ), .ZN(_05650_ ) );
AND3_X1 _13066_ ( .A1(_05609_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][10] ), .ZN(_05651_ ) );
AOI211_X1 _13067_ ( .A(fanout_net_10 ), .B(_05651_ ), .C1(\u_icache.cblocks[3][10] ), .C2(_05577_ ), .ZN(_05652_ ) );
OR2_X1 _13068_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][10] ), .ZN(_05653_ ) );
OR2_X1 _13069_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][10] ), .ZN(_05654_ ) );
NAND3_X1 _13070_ ( .A1(_05653_ ), .A2(_05511_ ), .A3(_05654_ ), .ZN(_05655_ ) );
AND3_X1 _13071_ ( .A1(_05559_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][10] ), .ZN(_05656_ ) );
AOI211_X1 _13072_ ( .A(_05625_ ), .B(_05656_ ), .C1(\u_icache.cblocks[7][10] ), .C2(_05604_ ), .ZN(_05657_ ) );
AOI221_X4 _13073_ ( .A(_05562_ ), .B1(_05650_ ), .B2(_05652_ ), .C1(_05655_ ), .C2(_05657_ ), .ZN(_00394_ ) );
OR2_X1 _13074_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][9] ), .ZN(_05658_ ) );
BUF_X4 _13075_ ( .A(_05484_ ), .Z(_05659_ ) );
OR2_X1 _13076_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][9] ), .ZN(_05660_ ) );
NAND3_X1 _13077_ ( .A1(_05658_ ), .A2(_05659_ ), .A3(_05660_ ), .ZN(_05661_ ) );
AND3_X1 _13078_ ( .A1(_05609_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][9] ), .ZN(_05662_ ) );
AOI211_X1 _13079_ ( .A(fanout_net_10 ), .B(_05662_ ), .C1(\u_icache.cblocks[3][9] ), .C2(_05577_ ), .ZN(_05663_ ) );
OR2_X1 _13080_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][9] ), .ZN(_05664_ ) );
OR2_X1 _13081_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][9] ), .ZN(_05665_ ) );
NAND3_X1 _13082_ ( .A1(_05664_ ), .A2(_05511_ ), .A3(_05665_ ), .ZN(_05666_ ) );
CLKBUF_X2 _13083_ ( .A(_05480_ ), .Z(_05667_ ) );
AND3_X1 _13084_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][9] ), .ZN(_05668_ ) );
AOI211_X1 _13085_ ( .A(_05625_ ), .B(_05668_ ), .C1(\u_icache.cblocks[7][9] ), .C2(_05604_ ), .ZN(_05669_ ) );
AOI221_X4 _13086_ ( .A(_05562_ ), .B1(_05661_ ), .B2(_05663_ ), .C1(_05666_ ), .C2(_05669_ ), .ZN(_00395_ ) );
BUF_X4 _13087_ ( .A(_05477_ ), .Z(_05670_ ) );
AND2_X1 _13088_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][8] ), .ZN(_05671_ ) );
AND2_X1 _13089_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[1][8] ), .ZN(_05672_ ) );
OAI21_X1 _13090_ ( .A(_05528_ ), .B1(_05671_ ), .B2(_05672_ ), .ZN(_05673_ ) );
AND3_X1 _13091_ ( .A1(_05609_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][8] ), .ZN(_05674_ ) );
AOI211_X1 _13092_ ( .A(fanout_net_10 ), .B(_05674_ ), .C1(\u_icache.cblocks[3][8] ), .C2(_05577_ ), .ZN(_05675_ ) );
OR2_X1 _13093_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][8] ), .ZN(_05676_ ) );
OR2_X1 _13094_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][8] ), .ZN(_05677_ ) );
NAND3_X1 _13095_ ( .A1(_05676_ ), .A2(_05494_ ), .A3(_05677_ ), .ZN(_05678_ ) );
AND3_X1 _13096_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][8] ), .ZN(_05679_ ) );
AOI211_X1 _13097_ ( .A(_05625_ ), .B(_05679_ ), .C1(\u_icache.cblocks[7][8] ), .C2(_05604_ ), .ZN(_05680_ ) );
AOI221_X4 _13098_ ( .A(_05670_ ), .B1(_05673_ ), .B2(_05675_ ), .C1(_05678_ ), .C2(_05680_ ), .ZN(_00396_ ) );
OR2_X1 _13099_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][7] ), .ZN(_05681_ ) );
OR2_X1 _13100_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][7] ), .ZN(_05682_ ) );
NAND3_X1 _13101_ ( .A1(_05681_ ), .A2(_05659_ ), .A3(_05682_ ), .ZN(_05683_ ) );
AND3_X1 _13102_ ( .A1(_05609_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][7] ), .ZN(_05684_ ) );
BUF_X4 _13103_ ( .A(_05490_ ), .Z(_05685_ ) );
AOI211_X1 _13104_ ( .A(fanout_net_10 ), .B(_05684_ ), .C1(\u_icache.cblocks[3][7] ), .C2(_05685_ ), .ZN(_05686_ ) );
OR2_X1 _13105_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][7] ), .ZN(_05687_ ) );
OR2_X1 _13106_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][7] ), .ZN(_05688_ ) );
NAND3_X1 _13107_ ( .A1(_05687_ ), .A2(_05494_ ), .A3(_05688_ ), .ZN(_05689_ ) );
AND3_X1 _13108_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][7] ), .ZN(_05690_ ) );
AOI211_X1 _13109_ ( .A(_05625_ ), .B(_05690_ ), .C1(\u_icache.cblocks[7][7] ), .C2(_05604_ ), .ZN(_05691_ ) );
AOI221_X4 _13110_ ( .A(_05670_ ), .B1(_05683_ ), .B2(_05686_ ), .C1(_05689_ ), .C2(_05691_ ), .ZN(_00397_ ) );
AND2_X1 _13111_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][6] ), .ZN(_05692_ ) );
AND2_X1 _13112_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[1][6] ), .ZN(_05693_ ) );
OAI21_X1 _13113_ ( .A(_05528_ ), .B1(_05692_ ), .B2(_05693_ ), .ZN(_05694_ ) );
AND3_X1 _13114_ ( .A1(_05609_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][6] ), .ZN(_05695_ ) );
AOI211_X1 _13115_ ( .A(fanout_net_10 ), .B(_05695_ ), .C1(\u_icache.cblocks[3][6] ), .C2(_05685_ ), .ZN(_05696_ ) );
AND2_X1 _13116_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][6] ), .ZN(_05697_ ) );
AND2_X1 _13117_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[5][6] ), .ZN(_05698_ ) );
OAI21_X1 _13118_ ( .A(_05545_ ), .B1(_05697_ ), .B2(_05698_ ), .ZN(_05699_ ) );
AND3_X1 _13119_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][6] ), .ZN(_05700_ ) );
AOI211_X1 _13120_ ( .A(_05625_ ), .B(_05700_ ), .C1(\u_icache.cblocks[7][6] ), .C2(_05604_ ), .ZN(_05701_ ) );
AOI221_X4 _13121_ ( .A(_05670_ ), .B1(_05694_ ), .B2(_05696_ ), .C1(_05699_ ), .C2(_05701_ ), .ZN(_00398_ ) );
OR2_X1 _13122_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][5] ), .ZN(_05702_ ) );
OR2_X1 _13123_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][5] ), .ZN(_05703_ ) );
NAND3_X1 _13124_ ( .A1(_05702_ ), .A2(_05659_ ), .A3(_05703_ ), .ZN(_05704_ ) );
AND3_X1 _13125_ ( .A1(_05609_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][5] ), .ZN(_05705_ ) );
AOI211_X1 _13126_ ( .A(fanout_net_10 ), .B(_05705_ ), .C1(\u_icache.cblocks[3][5] ), .C2(_05685_ ), .ZN(_05706_ ) );
AND2_X1 _13127_ ( .A1(_05496_ ), .A2(\u_icache.cblocks[4][5] ), .ZN(_05707_ ) );
AND2_X1 _13128_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[5][5] ), .ZN(_05708_ ) );
OAI21_X1 _13129_ ( .A(_05545_ ), .B1(_05707_ ), .B2(_05708_ ), .ZN(_05709_ ) );
AND3_X1 _13130_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][5] ), .ZN(_05710_ ) );
BUF_X4 _13131_ ( .A(_05491_ ), .Z(_05711_ ) );
AOI211_X1 _13132_ ( .A(_05625_ ), .B(_05710_ ), .C1(\u_icache.cblocks[7][5] ), .C2(_05711_ ), .ZN(_05712_ ) );
AOI221_X4 _13133_ ( .A(_05670_ ), .B1(_05704_ ), .B2(_05706_ ), .C1(_05709_ ), .C2(_05712_ ), .ZN(_00399_ ) );
OR2_X1 _13134_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][4] ), .ZN(_05713_ ) );
OR2_X1 _13135_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][4] ), .ZN(_05714_ ) );
NAND3_X1 _13136_ ( .A1(_05713_ ), .A2(_05659_ ), .A3(_05714_ ), .ZN(_05715_ ) );
CLKBUF_X2 _13137_ ( .A(_05479_ ), .Z(_05716_ ) );
AND3_X1 _13138_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][4] ), .ZN(_05717_ ) );
AOI211_X1 _13139_ ( .A(fanout_net_10 ), .B(_05717_ ), .C1(\u_icache.cblocks[3][4] ), .C2(_05685_ ), .ZN(_05718_ ) );
OR2_X1 _13140_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][4] ), .ZN(_05719_ ) );
OR2_X1 _13141_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][4] ), .ZN(_05720_ ) );
NAND3_X1 _13142_ ( .A1(_05719_ ), .A2(_05494_ ), .A3(_05720_ ), .ZN(_05721_ ) );
AND3_X1 _13143_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][4] ), .ZN(_05722_ ) );
AOI211_X1 _13144_ ( .A(_05625_ ), .B(_05722_ ), .C1(\u_icache.cblocks[7][4] ), .C2(_05711_ ), .ZN(_05723_ ) );
AOI221_X4 _13145_ ( .A(_05670_ ), .B1(_05715_ ), .B2(_05718_ ), .C1(_05721_ ), .C2(_05723_ ), .ZN(_00400_ ) );
AND2_X1 _13146_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][3] ), .ZN(_05724_ ) );
AND2_X1 _13147_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[1][3] ), .ZN(_05725_ ) );
OAI21_X1 _13148_ ( .A(_05484_ ), .B1(_05724_ ), .B2(_05725_ ), .ZN(_05726_ ) );
AND3_X1 _13149_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][3] ), .ZN(_05727_ ) );
AOI211_X1 _13150_ ( .A(fanout_net_10 ), .B(_05727_ ), .C1(\u_icache.cblocks[3][3] ), .C2(_05685_ ), .ZN(_05728_ ) );
AND2_X1 _13151_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[4][3] ), .ZN(_05729_ ) );
AND2_X1 _13152_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[5][3] ), .ZN(_05730_ ) );
OAI21_X1 _13153_ ( .A(_05545_ ), .B1(_05729_ ), .B2(_05730_ ), .ZN(_05731_ ) );
BUF_X4 _13154_ ( .A(_05468_ ), .Z(_05732_ ) );
AND3_X1 _13155_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][3] ), .ZN(_05733_ ) );
AOI211_X1 _13156_ ( .A(_05732_ ), .B(_05733_ ), .C1(\u_icache.cblocks[7][3] ), .C2(_05711_ ), .ZN(_05734_ ) );
AOI221_X4 _13157_ ( .A(_05670_ ), .B1(_05726_ ), .B2(_05728_ ), .C1(_05731_ ), .C2(_05734_ ), .ZN(_00401_ ) );
OR2_X1 _13158_ ( .A1(_05517_ ), .A2(\u_icache.cblocks[1][2] ), .ZN(_05735_ ) );
OR2_X1 _13159_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][2] ), .ZN(_05736_ ) );
NAND3_X1 _13160_ ( .A1(_05735_ ), .A2(_05659_ ), .A3(_05736_ ), .ZN(_05737_ ) );
AND3_X1 _13161_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][2] ), .ZN(_05738_ ) );
AOI211_X1 _13162_ ( .A(fanout_net_10 ), .B(_05738_ ), .C1(\u_icache.cblocks[3][2] ), .C2(_05685_ ), .ZN(_05739_ ) );
AND2_X1 _13163_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[4][2] ), .ZN(_05740_ ) );
AND2_X1 _13164_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[5][2] ), .ZN(_05741_ ) );
OAI21_X1 _13165_ ( .A(_05545_ ), .B1(_05740_ ), .B2(_05741_ ), .ZN(_05742_ ) );
AND3_X1 _13166_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][2] ), .ZN(_05743_ ) );
AOI211_X1 _13167_ ( .A(_05732_ ), .B(_05743_ ), .C1(\u_icache.cblocks[7][2] ), .C2(_05711_ ), .ZN(_05744_ ) );
AOI221_X4 _13168_ ( .A(_05670_ ), .B1(_05737_ ), .B2(_05739_ ), .C1(_05742_ ), .C2(_05744_ ), .ZN(_00402_ ) );
OR2_X1 _13169_ ( .A1(_05500_ ), .A2(\u_icache.cblocks[1][28] ), .ZN(_05745_ ) );
OR2_X1 _13170_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][28] ), .ZN(_05746_ ) );
NAND3_X1 _13171_ ( .A1(_05745_ ), .A2(_05659_ ), .A3(_05746_ ), .ZN(_05747_ ) );
AND3_X1 _13172_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][28] ), .ZN(_05748_ ) );
AOI211_X1 _13173_ ( .A(fanout_net_10 ), .B(_05748_ ), .C1(\u_icache.cblocks[3][28] ), .C2(_05685_ ), .ZN(_05749_ ) );
OR2_X1 _13174_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][28] ), .ZN(_05750_ ) );
OR2_X1 _13175_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][28] ), .ZN(_05751_ ) );
NAND3_X1 _13176_ ( .A1(_05750_ ), .A2(_05494_ ), .A3(_05751_ ), .ZN(_05752_ ) );
AND3_X1 _13177_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][28] ), .ZN(_05753_ ) );
AOI211_X1 _13178_ ( .A(_05732_ ), .B(_05753_ ), .C1(\u_icache.cblocks[7][28] ), .C2(_05711_ ), .ZN(_05754_ ) );
AOI221_X4 _13179_ ( .A(_05670_ ), .B1(_05747_ ), .B2(_05749_ ), .C1(_05752_ ), .C2(_05754_ ), .ZN(_00403_ ) );
OR2_X1 _13180_ ( .A1(_05500_ ), .A2(\u_icache.cblocks[1][1] ), .ZN(_05755_ ) );
OR2_X1 _13181_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][1] ), .ZN(_05756_ ) );
NAND3_X1 _13182_ ( .A1(_05755_ ), .A2(_05659_ ), .A3(_05756_ ), .ZN(_05757_ ) );
AND3_X1 _13183_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][1] ), .ZN(_05758_ ) );
AOI211_X1 _13184_ ( .A(fanout_net_10 ), .B(_05758_ ), .C1(\u_icache.cblocks[3][1] ), .C2(_05685_ ), .ZN(_05759_ ) );
OR2_X1 _13185_ ( .A1(_05599_ ), .A2(\u_icache.cblocks[5][1] ), .ZN(_05760_ ) );
OR2_X1 _13186_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][1] ), .ZN(_05761_ ) );
NAND3_X1 _13187_ ( .A1(_05760_ ), .A2(_05494_ ), .A3(_05761_ ), .ZN(_05762_ ) );
AND3_X1 _13188_ ( .A1(_05667_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][1] ), .ZN(_05763_ ) );
AOI211_X1 _13189_ ( .A(_05732_ ), .B(_05763_ ), .C1(\u_icache.cblocks[7][1] ), .C2(_05711_ ), .ZN(_05764_ ) );
AOI221_X4 _13190_ ( .A(_05670_ ), .B1(_05757_ ), .B2(_05759_ ), .C1(_05762_ ), .C2(_05764_ ), .ZN(_00404_ ) );
AND2_X1 _13191_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][0] ), .ZN(_05765_ ) );
AND2_X1 _13192_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[1][0] ), .ZN(_05766_ ) );
OAI21_X1 _13193_ ( .A(_05484_ ), .B1(_05765_ ), .B2(_05766_ ), .ZN(_05767_ ) );
AND3_X1 _13194_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][0] ), .ZN(_05768_ ) );
AOI211_X1 _13195_ ( .A(fanout_net_10 ), .B(_05768_ ), .C1(\u_icache.cblocks[3][0] ), .C2(_05685_ ), .ZN(_05769_ ) );
OR2_X1 _13196_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[5][0] ), .ZN(_05770_ ) );
OR2_X1 _13197_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][0] ), .ZN(_05771_ ) );
NAND3_X1 _13198_ ( .A1(_05770_ ), .A2(_05494_ ), .A3(_05771_ ), .ZN(_05772_ ) );
AND3_X1 _13199_ ( .A1(_05495_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][0] ), .ZN(_05773_ ) );
AOI211_X1 _13200_ ( .A(_05732_ ), .B(_05773_ ), .C1(\u_icache.cblocks[7][0] ), .C2(_05711_ ), .ZN(_05774_ ) );
AOI221_X4 _13201_ ( .A(_05670_ ), .B1(_05767_ ), .B2(_05769_ ), .C1(_05772_ ), .C2(_05774_ ), .ZN(_00405_ ) );
AND2_X1 _13202_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][27] ), .ZN(_05775_ ) );
AND2_X1 _13203_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[1][27] ), .ZN(_05776_ ) );
OAI21_X1 _13204_ ( .A(_05484_ ), .B1(_05775_ ), .B2(_05776_ ), .ZN(_05777_ ) );
AND3_X1 _13205_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][27] ), .ZN(_05778_ ) );
AOI211_X1 _13206_ ( .A(fanout_net_10 ), .B(_05778_ ), .C1(\u_icache.cblocks[3][27] ), .C2(_05685_ ), .ZN(_05779_ ) );
AND2_X1 _13207_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[4][27] ), .ZN(_05780_ ) );
AND2_X1 _13208_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[5][27] ), .ZN(_05781_ ) );
OAI21_X1 _13209_ ( .A(_05545_ ), .B1(_05780_ ), .B2(_05781_ ), .ZN(_05782_ ) );
AND3_X1 _13210_ ( .A1(_05495_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][27] ), .ZN(_05783_ ) );
AOI211_X1 _13211_ ( .A(_05732_ ), .B(_05783_ ), .C1(\u_icache.cblocks[7][27] ), .C2(_05711_ ), .ZN(_05784_ ) );
AOI221_X4 _13212_ ( .A(_05477_ ), .B1(_05777_ ), .B2(_05779_ ), .C1(_05782_ ), .C2(_05784_ ), .ZN(_00406_ ) );
OR2_X1 _13213_ ( .A1(_05500_ ), .A2(\u_icache.cblocks[1][26] ), .ZN(_05785_ ) );
OR2_X1 _13214_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][26] ), .ZN(_05786_ ) );
NAND3_X1 _13215_ ( .A1(_05785_ ), .A2(_05659_ ), .A3(_05786_ ), .ZN(_05787_ ) );
AND3_X1 _13216_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][26] ), .ZN(_05788_ ) );
AOI211_X1 _13217_ ( .A(fanout_net_10 ), .B(_05788_ ), .C1(\u_icache.cblocks[3][26] ), .C2(_05491_ ), .ZN(_05789_ ) );
OR2_X1 _13218_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[5][26] ), .ZN(_05790_ ) );
OR2_X1 _13219_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][26] ), .ZN(_05791_ ) );
NAND3_X1 _13220_ ( .A1(_05790_ ), .A2(_05494_ ), .A3(_05791_ ), .ZN(_05792_ ) );
AND3_X1 _13221_ ( .A1(_05495_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][26] ), .ZN(_05793_ ) );
AOI211_X1 _13222_ ( .A(_05732_ ), .B(_05793_ ), .C1(\u_icache.cblocks[7][26] ), .C2(_05711_ ), .ZN(_05794_ ) );
AOI221_X4 _13223_ ( .A(_05477_ ), .B1(_05787_ ), .B2(_05789_ ), .C1(_05792_ ), .C2(_05794_ ), .ZN(_00407_ ) );
OR2_X1 _13224_ ( .A1(_05500_ ), .A2(\u_icache.cblocks[1][25] ), .ZN(_05795_ ) );
OR2_X1 _13225_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[0][25] ), .ZN(_05796_ ) );
NAND3_X1 _13226_ ( .A1(_05795_ ), .A2(_05659_ ), .A3(_05796_ ), .ZN(_05797_ ) );
AND3_X1 _13227_ ( .A1(_05716_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[2][25] ), .ZN(_05798_ ) );
AOI211_X1 _13228_ ( .A(fanout_net_10 ), .B(_05798_ ), .C1(\u_icache.cblocks[3][25] ), .C2(_05491_ ), .ZN(_05799_ ) );
OR2_X1 _13229_ ( .A1(_05529_ ), .A2(\u_icache.cblocks[5][25] ), .ZN(_05800_ ) );
OR2_X1 _13230_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][25] ), .ZN(_05801_ ) );
NAND3_X1 _13231_ ( .A1(_05800_ ), .A2(_05494_ ), .A3(_05801_ ), .ZN(_05802_ ) );
AND3_X1 _13232_ ( .A1(_05495_ ), .A2(fanout_net_9 ), .A3(\u_icache.cblocks[6][25] ), .ZN(_05803_ ) );
AOI211_X1 _13233_ ( .A(_05732_ ), .B(_05803_ ), .C1(\u_icache.cblocks[7][25] ), .C2(_05711_ ), .ZN(_05804_ ) );
AOI221_X4 _13234_ ( .A(_05477_ ), .B1(_05797_ ), .B2(_05799_ ), .C1(_05802_ ), .C2(_05804_ ), .ZN(_00408_ ) );
OR2_X1 _13235_ ( .A1(_05500_ ), .A2(\u_icache.cblocks[1][24] ), .ZN(_05805_ ) );
OR2_X1 _13236_ ( .A1(\fc_addr[2] ), .A2(\u_icache.cblocks[0][24] ), .ZN(_05806_ ) );
NAND3_X1 _13237_ ( .A1(_05805_ ), .A2(_05659_ ), .A3(_05806_ ), .ZN(_05807_ ) );
AND3_X1 _13238_ ( .A1(_05716_ ), .A2(\fc_addr[3] ), .A3(\u_icache.cblocks[2][24] ), .ZN(_05808_ ) );
AOI211_X1 _13239_ ( .A(\fc_addr[4] ), .B(_05808_ ), .C1(\u_icache.cblocks[3][24] ), .C2(_05491_ ), .ZN(_05809_ ) );
AND2_X1 _13240_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[4][24] ), .ZN(_05810_ ) );
AND2_X1 _13241_ ( .A1(\fc_addr[2] ), .A2(\u_icache.cblocks[5][24] ), .ZN(_05811_ ) );
OAI21_X1 _13242_ ( .A(_05485_ ), .B1(_05810_ ), .B2(_05811_ ), .ZN(_05812_ ) );
AND3_X1 _13243_ ( .A1(_05495_ ), .A2(\fc_addr[3] ), .A3(\u_icache.cblocks[6][24] ), .ZN(_05813_ ) );
AOI211_X1 _13244_ ( .A(_05732_ ), .B(_05813_ ), .C1(\u_icache.cblocks[7][24] ), .C2(_05492_ ), .ZN(_05814_ ) );
AOI221_X4 _13245_ ( .A(_05477_ ), .B1(_05807_ ), .B2(_05809_ ), .C1(_05812_ ), .C2(_05814_ ), .ZN(_00409_ ) );
AND2_X1 _13246_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][23] ), .ZN(_05815_ ) );
AND2_X1 _13247_ ( .A1(\fc_addr[2] ), .A2(\u_icache.cblocks[1][23] ), .ZN(_05816_ ) );
OAI21_X1 _13248_ ( .A(_05484_ ), .B1(_05815_ ), .B2(_05816_ ), .ZN(_05817_ ) );
AND3_X1 _13249_ ( .A1(_05480_ ), .A2(\fc_addr[3] ), .A3(\u_icache.cblocks[2][23] ), .ZN(_05818_ ) );
AOI211_X1 _13250_ ( .A(\fc_addr[4] ), .B(_05818_ ), .C1(\u_icache.cblocks[3][23] ), .C2(_05491_ ), .ZN(_05819_ ) );
AND2_X1 _13251_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[4][23] ), .ZN(_05820_ ) );
AND2_X1 _13252_ ( .A1(\fc_addr[2] ), .A2(\u_icache.cblocks[5][23] ), .ZN(_05821_ ) );
OAI21_X1 _13253_ ( .A(_05485_ ), .B1(_05820_ ), .B2(_05821_ ), .ZN(_05822_ ) );
AND3_X1 _13254_ ( .A1(_05495_ ), .A2(\fc_addr[3] ), .A3(\u_icache.cblocks[6][23] ), .ZN(_05823_ ) );
AOI211_X1 _13255_ ( .A(_05732_ ), .B(_05823_ ), .C1(\u_icache.cblocks[7][23] ), .C2(_05492_ ), .ZN(_05824_ ) );
AOI221_X4 _13256_ ( .A(_05477_ ), .B1(_05817_ ), .B2(_05819_ ), .C1(_05822_ ), .C2(_05824_ ), .ZN(_00410_ ) );
AND2_X1 _13257_ ( .A1(_05481_ ), .A2(\u_icache.cblocks[0][22] ), .ZN(_05825_ ) );
AND2_X1 _13258_ ( .A1(\fc_addr[2] ), .A2(\u_icache.cblocks[1][22] ), .ZN(_05826_ ) );
OAI21_X1 _13259_ ( .A(_05484_ ), .B1(_05825_ ), .B2(_05826_ ), .ZN(_05827_ ) );
AND3_X1 _13260_ ( .A1(_05480_ ), .A2(\fc_addr[3] ), .A3(\u_icache.cblocks[2][22] ), .ZN(_05828_ ) );
AOI211_X1 _13261_ ( .A(\fc_addr[4] ), .B(_05828_ ), .C1(\u_icache.cblocks[3][22] ), .C2(_05491_ ), .ZN(_05829_ ) );
AND2_X1 _13262_ ( .A1(_05509_ ), .A2(\u_icache.cblocks[4][22] ), .ZN(_05830_ ) );
AND2_X1 _13263_ ( .A1(\fc_addr[2] ), .A2(\u_icache.cblocks[5][22] ), .ZN(_05831_ ) );
OAI21_X1 _13264_ ( .A(_05485_ ), .B1(_05830_ ), .B2(_05831_ ), .ZN(_05832_ ) );
AND3_X1 _13265_ ( .A1(_05495_ ), .A2(\fc_addr[3] ), .A3(\u_icache.cblocks[6][22] ), .ZN(_05833_ ) );
AOI211_X1 _13266_ ( .A(_05468_ ), .B(_05833_ ), .C1(\u_icache.cblocks[7][22] ), .C2(_05492_ ), .ZN(_05834_ ) );
AOI221_X4 _13267_ ( .A(_05477_ ), .B1(_05827_ ), .B2(_05829_ ), .C1(_05832_ ), .C2(_05834_ ), .ZN(_00411_ ) );
INV_X1 _13268_ ( .A(_00760_ ), .ZN(_05835_ ) );
OAI21_X1 _13269_ ( .A(\u_ifu.jpc_ok_$_NOT__A_Y ), .B1(_05835_ ), .B2(_00742_ ), .ZN(_05836_ ) );
NAND4_X1 _13270_ ( .A1(_00745_ ), .A2(idu_ready ), .A3(_00761_ ), .A4(_00759_ ), .ZN(_05837_ ) );
INV_X1 _13271_ ( .A(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ), .ZN(_05838_ ) );
INV_X1 _13272_ ( .A(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .ZN(_05839_ ) );
NAND2_X1 _13273_ ( .A1(_05839_ ), .A2(\u_icache.ctags[0][5] ), .ZN(_05840_ ) );
NAND2_X1 _13274_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][5] ), .ZN(_05841_ ) );
AND3_X1 _13275_ ( .A1(_05840_ ), .A2(\fc_addr[10] ), .A3(_05841_ ), .ZN(_05842_ ) );
MUX2_X1 _13276_ ( .A(\u_icache.ctags[0][16] ), .B(\u_icache.ctags[1][16] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05843_ ) );
AND2_X1 _13277_ ( .A1(_05843_ ), .A2(_05449_ ), .ZN(_05844_ ) );
MUX2_X1 _13278_ ( .A(\u_icache.ctags[0][10] ), .B(\u_icache.ctags[1][10] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05845_ ) );
NOR2_X1 _13279_ ( .A1(_05845_ ), .A2(_05455_ ), .ZN(_05846_ ) );
AOI21_X1 _13280_ ( .A(\fc_addr[10] ), .B1(_05840_ ), .B2(_05841_ ), .ZN(_05847_ ) );
OR4_X1 _13281_ ( .A1(_05842_ ), .A2(_05844_ ), .A3(_05846_ ), .A4(_05847_ ), .ZN(_05848_ ) );
MUX2_X1 _13282_ ( .A(\u_icache.ctags[0][19] ), .B(\u_icache.ctags[1][19] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05849_ ) );
MUX2_X1 _13283_ ( .A(\u_icache.ctags[0][17] ), .B(\u_icache.ctags[1][17] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05850_ ) );
AOI22_X1 _13284_ ( .A1(_05474_ ), .A2(_05849_ ), .B1(_05850_ ), .B2(_05476_ ), .ZN(_05851_ ) );
MUX2_X1 _13285_ ( .A(\u_icache.ctags[0][23] ), .B(\u_icache.ctags[1][23] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05852_ ) );
INV_X1 _13286_ ( .A(_05852_ ), .ZN(_05853_ ) );
OAI221_X1 _13287_ ( .A(_05851_ ), .B1(\fc_addr[28] ), .B2(_05853_ ), .C1(_05476_ ), .C2(_05850_ ), .ZN(_05854_ ) );
NOR2_X1 _13288_ ( .A1(_05848_ ), .A2(_05854_ ), .ZN(_05855_ ) );
NAND2_X1 _13289_ ( .A1(_05839_ ), .A2(\u_icache.ctags[0][24] ), .ZN(_05856_ ) );
NAND2_X1 _13290_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][24] ), .ZN(_05857_ ) );
NAND2_X1 _13291_ ( .A1(_05856_ ), .A2(_05857_ ), .ZN(_05858_ ) );
AOI22_X1 _13292_ ( .A1(_05853_ ), .A2(\fc_addr[28] ), .B1(_05460_ ), .B2(_05858_ ), .ZN(_05859_ ) );
MUX2_X1 _13293_ ( .A(\u_icache.ctags[0][25] ), .B(\u_icache.ctags[1][25] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05860_ ) );
MUX2_X1 _13294_ ( .A(\u_icache.ctags[0][12] ), .B(\u_icache.ctags[1][12] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05861_ ) );
OAI221_X1 _13295_ ( .A(_05859_ ), .B1(_05448_ ), .B2(_05860_ ), .C1(_05453_ ), .C2(_05861_ ), .ZN(_05862_ ) );
AND2_X1 _13296_ ( .A1(_05845_ ), .A2(_05455_ ), .ZN(_05863_ ) );
NOR2_X1 _13297_ ( .A1(_05849_ ), .A2(_05474_ ), .ZN(_05864_ ) );
NAND2_X1 _13298_ ( .A1(_05839_ ), .A2(\u_icache.ctags[0][9] ), .ZN(_05865_ ) );
NAND2_X1 _13299_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][9] ), .ZN(_05866_ ) );
AND3_X1 _13300_ ( .A1(_05865_ ), .A2(\fc_addr[14] ), .A3(_05866_ ), .ZN(_05867_ ) );
AOI21_X1 _13301_ ( .A(\fc_addr[14] ), .B1(_05865_ ), .B2(_05866_ ), .ZN(_05868_ ) );
OR4_X1 _13302_ ( .A1(_05863_ ), .A2(_05864_ ), .A3(_05867_ ), .A4(_05868_ ), .ZN(_05869_ ) );
MUX2_X1 _13303_ ( .A(\u_icache.ctags[0][14] ), .B(\u_icache.ctags[1][14] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05870_ ) );
AOI22_X1 _13304_ ( .A1(_05451_ ), .A2(_05870_ ), .B1(_05861_ ), .B2(_05453_ ), .ZN(_05871_ ) );
MUX2_X1 _13305_ ( .A(\u_icache.ctags[0][4] ), .B(\u_icache.ctags[1][4] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05872_ ) );
OAI221_X1 _13306_ ( .A(_05871_ ), .B1(_05449_ ), .B2(_05843_ ), .C1(_05463_ ), .C2(_05872_ ), .ZN(_05873_ ) );
MUX2_X1 _13307_ ( .A(\u_icache.ctags[0][8] ), .B(\u_icache.ctags[1][8] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05874_ ) );
MUX2_X1 _13308_ ( .A(\u_icache.ctags[0][21] ), .B(\u_icache.ctags[1][21] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05875_ ) );
AOI22_X1 _13309_ ( .A1(_05458_ ), .A2(_05874_ ), .B1(_05875_ ), .B2(_05472_ ), .ZN(_05876_ ) );
OR2_X1 _13310_ ( .A1(_05874_ ), .A2(_05458_ ), .ZN(_05877_ ) );
OAI211_X1 _13311_ ( .A(_05876_ ), .B(_05877_ ), .C1(_05472_ ), .C2(_05875_ ), .ZN(_05878_ ) );
NOR4_X1 _13312_ ( .A1(_05862_ ), .A2(_05869_ ), .A3(_05873_ ), .A4(_05878_ ), .ZN(_05879_ ) );
BUF_X4 _13313_ ( .A(_05839_ ), .Z(_05880_ ) );
NAND2_X1 _13314_ ( .A1(_05880_ ), .A2(\u_icache.ctags[0][18] ), .ZN(_05881_ ) );
NAND2_X1 _13315_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][18] ), .ZN(_05882_ ) );
AND3_X1 _13316_ ( .A1(_05881_ ), .A2(\fc_addr[23] ), .A3(_05882_ ), .ZN(_05883_ ) );
AOI21_X1 _13317_ ( .A(\fc_addr[23] ), .B1(_05881_ ), .B2(_05882_ ), .ZN(_05884_ ) );
NAND2_X1 _13318_ ( .A1(_05880_ ), .A2(\u_icache.ctags[0][20] ), .ZN(_05885_ ) );
NAND2_X1 _13319_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][20] ), .ZN(_05886_ ) );
AOI21_X1 _13320_ ( .A(\fc_addr[25] ), .B1(_05885_ ), .B2(_05886_ ), .ZN(_05887_ ) );
NOR3_X1 _13321_ ( .A1(_05883_ ), .A2(_05884_ ), .A3(_05887_ ), .ZN(_05888_ ) );
AND3_X1 _13322_ ( .A1(_05885_ ), .A2(\fc_addr[25] ), .A3(_05886_ ), .ZN(_05889_ ) );
NAND2_X1 _13323_ ( .A1(_05839_ ), .A2(\u_icache.ctags[0][15] ), .ZN(_05890_ ) );
NAND2_X1 _13324_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][15] ), .ZN(_05891_ ) );
NAND2_X1 _13325_ ( .A1(_05890_ ), .A2(_05891_ ), .ZN(_05892_ ) );
XNOR2_X1 _13326_ ( .A(_05892_ ), .B(_05450_ ), .ZN(_05893_ ) );
AOI211_X1 _13327_ ( .A(_05889_ ), .B(_05893_ ), .C1(_05448_ ), .C2(_05860_ ), .ZN(_05894_ ) );
AND4_X1 _13328_ ( .A1(_05855_ ), .A2(_05879_ ), .A3(_05888_ ), .A4(_05894_ ), .ZN(_05895_ ) );
MUX2_X1 _13329_ ( .A(\u_icache.ctags[0][1] ), .B(\u_icache.ctags[1][1] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05896_ ) );
NOR2_X1 _13330_ ( .A1(_05896_ ), .A2(_05466_ ), .ZN(_05897_ ) );
AOI21_X1 _13331_ ( .A(_05897_ ), .B1(_05463_ ), .B2(_05872_ ), .ZN(_05898_ ) );
MUX2_X1 _13332_ ( .A(\u_icache.ctags[0][6] ), .B(\u_icache.ctags[1][6] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05899_ ) );
NAND2_X1 _13333_ ( .A1(_05899_ ), .A2(_05461_ ), .ZN(_05900_ ) );
OAI211_X1 _13334_ ( .A(_05898_ ), .B(_05900_ ), .C1(_05460_ ), .C2(_05858_ ), .ZN(_05901_ ) );
NOR2_X1 _13335_ ( .A1(_05880_ ), .A2(\u_icache.ctags[1][3] ), .ZN(_05902_ ) );
NOR2_X1 _13336_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[0][3] ), .ZN(_05903_ ) );
NOR2_X1 _13337_ ( .A1(_05902_ ), .A2(_05903_ ), .ZN(_05904_ ) );
XNOR2_X1 _13338_ ( .A(_05904_ ), .B(\fc_addr[8] ), .ZN(_05905_ ) );
NOR2_X1 _13339_ ( .A1(_05880_ ), .A2(\u_icache.ctags[1][7] ), .ZN(_05906_ ) );
NOR2_X1 _13340_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[0][7] ), .ZN(_05907_ ) );
NOR2_X1 _13341_ ( .A1(_05906_ ), .A2(_05907_ ), .ZN(_05908_ ) );
XNOR2_X1 _13342_ ( .A(_05908_ ), .B(\fc_addr[12] ), .ZN(_05909_ ) );
NOR2_X1 _13343_ ( .A1(_05880_ ), .A2(\u_icache.ctags[1][11] ), .ZN(_05910_ ) );
NOR2_X1 _13344_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[0][11] ), .ZN(_05911_ ) );
NOR2_X1 _13345_ ( .A1(_05910_ ), .A2(_05911_ ), .ZN(_05912_ ) );
XNOR2_X1 _13346_ ( .A(_05912_ ), .B(\fc_addr[16] ), .ZN(_05913_ ) );
NAND2_X1 _13347_ ( .A1(_05880_ ), .A2(\u_icache.ctags[0][26] ), .ZN(_05914_ ) );
NAND2_X1 _13348_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][26] ), .ZN(_05915_ ) );
NAND2_X1 _13349_ ( .A1(_05914_ ), .A2(_05915_ ), .ZN(_05916_ ) );
XNOR2_X1 _13350_ ( .A(_05916_ ), .B(\fc_addr[31] ), .ZN(_05917_ ) );
NAND4_X1 _13351_ ( .A1(_05905_ ), .A2(_05909_ ), .A3(_05913_ ), .A4(_05917_ ), .ZN(_05918_ ) );
NOR2_X1 _13352_ ( .A1(_05880_ ), .A2(\u_icache.ctags[1][2] ), .ZN(_05919_ ) );
NOR2_X1 _13353_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[0][2] ), .ZN(_05920_ ) );
NOR2_X1 _13354_ ( .A1(_05919_ ), .A2(_05920_ ), .ZN(_05921_ ) );
XNOR2_X1 _13355_ ( .A(_05921_ ), .B(\fc_addr[7] ), .ZN(_05922_ ) );
NOR2_X1 _13356_ ( .A1(_05880_ ), .A2(\u_icache.ctags[1][22] ), .ZN(_05923_ ) );
NOR2_X1 _13357_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[0][22] ), .ZN(_05924_ ) );
NOR2_X1 _13358_ ( .A1(_05923_ ), .A2(_05924_ ), .ZN(_05925_ ) );
XNOR2_X1 _13359_ ( .A(_05925_ ), .B(\fc_addr[27] ), .ZN(_05926_ ) );
NAND2_X1 _13360_ ( .A1(_05880_ ), .A2(\u_icache.ctags[0][0] ), .ZN(_05927_ ) );
NAND2_X1 _13361_ ( .A1(\u_icache.ctags[1][0] ), .A2(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .ZN(_05928_ ) );
NAND2_X1 _13362_ ( .A1(_05927_ ), .A2(_05928_ ), .ZN(_05929_ ) );
XNOR2_X1 _13363_ ( .A(_05929_ ), .B(\fc_addr[5] ), .ZN(_05930_ ) );
NAND2_X1 _13364_ ( .A1(_05880_ ), .A2(\u_icache.ctags[0][13] ), .ZN(_05931_ ) );
NAND2_X1 _13365_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][13] ), .ZN(_05932_ ) );
NAND2_X1 _13366_ ( .A1(_05931_ ), .A2(_05932_ ), .ZN(_05933_ ) );
XNOR2_X1 _13367_ ( .A(_05933_ ), .B(\fc_addr[18] ), .ZN(_05934_ ) );
NAND4_X1 _13368_ ( .A1(_05922_ ), .A2(_05926_ ), .A3(_05930_ ), .A4(_05934_ ), .ZN(_05935_ ) );
OR2_X1 _13369_ ( .A1(_05899_ ), .A2(_05461_ ), .ZN(_05936_ ) );
OR2_X1 _13370_ ( .A1(_05870_ ), .A2(_05451_ ), .ZN(_05937_ ) );
MUX2_X1 _13371_ ( .A(\u_icache.cvalids[0] ), .B(\u_icache.cvalids[1] ), .S(\fc_addr[4] ), .Z(_05938_ ) );
NAND2_X1 _13372_ ( .A1(_05896_ ), .A2(_05466_ ), .ZN(_05939_ ) );
NAND4_X1 _13373_ ( .A1(_05936_ ), .A2(_05937_ ), .A3(_05938_ ), .A4(_05939_ ), .ZN(_05940_ ) );
NOR4_X1 _13374_ ( .A1(_05901_ ), .A2(_05918_ ), .A3(_05935_ ), .A4(_05940_ ), .ZN(_05941_ ) );
AOI211_X1 _13375_ ( .A(\u_icache.ended ), .B(_05838_ ), .C1(_05895_ ), .C2(_05941_ ), .ZN(_05942_ ) );
AND3_X1 _13376_ ( .A1(_05836_ ), .A2(_05837_ ), .A3(_05942_ ), .ZN(\u_icache.ended_$_ANDNOT__B_Y ) );
CLKBUF_X2 _13377_ ( .A(_00863_ ), .Z(_05943_ ) );
AND4_X1 _13378_ ( .A1(_05943_ ), .A2(_05836_ ), .A3(_05837_ ), .A4(_05942_ ), .ZN(_00412_ ) );
NOR2_X1 _13379_ ( .A1(_01215_ ), .A2(_01216_ ), .ZN(_05944_ ) );
AND2_X1 _13380_ ( .A1(\u_icache.count[1] ), .A2(\u_icache.count[0] ), .ZN(_05945_ ) );
INV_X1 _13381_ ( .A(\u_icache.count[2] ), .ZN(_05946_ ) );
XNOR2_X1 _13382_ ( .A(_05945_ ), .B(_05946_ ), .ZN(_05947_ ) );
AND4_X1 _13383_ ( .A1(_05943_ ), .A2(_05944_ ), .A3(_01195_ ), .A4(_05947_ ), .ZN(_00413_ ) );
AND2_X1 _13384_ ( .A1(_05944_ ), .A2(_01195_ ), .ZN(_05948_ ) );
INV_X1 _13385_ ( .A(_05948_ ), .ZN(_05949_ ) );
NOR2_X1 _13386_ ( .A1(\u_icache.count[1] ), .A2(\u_icache.count[0] ), .ZN(_05950_ ) );
NOR4_X1 _13387_ ( .A1(_05949_ ), .A2(_05478_ ), .A3(_05945_ ), .A4(_05950_ ), .ZN(_00414_ ) );
INV_X1 _13388_ ( .A(_05944_ ), .ZN(_05951_ ) );
NOR4_X1 _13389_ ( .A1(_05951_ ), .A2(\u_icache.count[0] ), .A3(_05478_ ), .A4(_01205_ ), .ZN(_00415_ ) );
INV_X1 _13390_ ( .A(ifu_ready ), .ZN(_05952_ ) );
AND3_X1 _13391_ ( .A1(_05895_ ), .A2(_05952_ ), .A3(_05941_ ), .ZN(_05953_ ) );
NAND3_X1 _13392_ ( .A1(_05836_ ), .A2(_05837_ ), .A3(_05953_ ), .ZN(_05954_ ) );
AND2_X1 _13393_ ( .A1(_05950_ ), .A2(\u_icache.count[2] ), .ZN(\u_icache.cvalids_$_SDFFE_PP0P__Q_E ) );
INV_X1 _13394_ ( .A(\u_icache.cvalids_$_SDFFE_PP0P__Q_E ), .ZN(_05955_ ) );
NAND2_X1 _13395_ ( .A1(_05954_ ), .A2(_05955_ ), .ZN(\u_icache.cready_$_ANDNOT__B_Y_$_OR__B_Y ) );
AOI21_X1 _13396_ ( .A(_04454_ ), .B1(_05954_ ), .B2(_05955_ ), .ZN(_00416_ ) );
NAND2_X1 _13397_ ( .A1(_05943_ ), .A2(\u_icache.cvalids[1] ), .ZN(_05956_ ) );
OAI21_X1 _13398_ ( .A(_05956_ ), .B1(_05478_ ), .B2(_05469_ ), .ZN(_00417_ ) );
NOR2_X1 _13399_ ( .A1(_05469_ ), .A2(\u_icache.cvalids[0] ), .ZN(_05957_ ) );
NOR3_X1 _13400_ ( .A1(_00857_ ), .A2(fanout_net_3 ), .A3(_05957_ ), .ZN(_00418_ ) );
AND4_X1 _13401_ ( .A1(_05946_ ), .A2(_05948_ ), .A3(_01060_ ), .A4(_05945_ ), .ZN(_00419_ ) );
BUF_X2 _13402_ ( .A(_00771_ ), .Z(\u_ifu.inst_ok_$_ANDNOT__A_Y ) );
INV_X1 _13403_ ( .A(_00770_ ), .ZN(_05958_ ) );
BUF_X4 _13404_ ( .A(_05958_ ), .Z(_05959_ ) );
NOR4_X1 _13405_ ( .A1(_04463_ ), .A2(fanout_net_3 ), .A3(_04462_ ), .A4(_05959_ ), .ZN(_00420_ ) );
AND3_X1 _13406_ ( .A1(_04461_ ), .A2(\fd_inst[31] ), .A3(_04464_ ), .ZN(_00421_ ) );
AND3_X1 _13407_ ( .A1(_04461_ ), .A2(\fd_inst[30] ), .A3(_04464_ ), .ZN(_00422_ ) );
CLKBUF_X2 _13408_ ( .A(_00864_ ), .Z(_05960_ ) );
AND3_X1 _13409_ ( .A1(_05960_ ), .A2(\fd_inst[21] ), .A3(_04464_ ), .ZN(_00423_ ) );
AND3_X1 _13410_ ( .A1(_05960_ ), .A2(\fd_inst[20] ), .A3(_04464_ ), .ZN(_00424_ ) );
AND3_X1 _13411_ ( .A1(_05960_ ), .A2(\fd_inst[19] ), .A3(_04464_ ), .ZN(_00425_ ) );
AND3_X1 _13412_ ( .A1(_05960_ ), .A2(\fd_inst[18] ), .A3(_04464_ ), .ZN(_00426_ ) );
AND3_X1 _13413_ ( .A1(_05960_ ), .A2(\fd_inst[17] ), .A3(_04464_ ), .ZN(_00427_ ) );
AND3_X1 _13414_ ( .A1(_05960_ ), .A2(\fd_inst[16] ), .A3(_04464_ ), .ZN(_00428_ ) );
CLKBUF_X2 _13415_ ( .A(_00637_ ), .Z(_05961_ ) );
AND3_X1 _13416_ ( .A1(_05960_ ), .A2(\fd_inst[15] ), .A3(_05961_ ), .ZN(_00429_ ) );
AND3_X1 _13417_ ( .A1(_05960_ ), .A2(\fd_inst[14] ), .A3(_05961_ ), .ZN(_00430_ ) );
AND3_X1 _13418_ ( .A1(_05960_ ), .A2(\fd_inst[13] ), .A3(_05961_ ), .ZN(_00431_ ) );
AND3_X1 _13419_ ( .A1(_05960_ ), .A2(\fd_inst[12] ), .A3(_05961_ ), .ZN(_00432_ ) );
CLKBUF_X2 _13420_ ( .A(_00864_ ), .Z(_05962_ ) );
AND3_X1 _13421_ ( .A1(_05962_ ), .A2(\fd_inst[29] ), .A3(_05961_ ), .ZN(_00433_ ) );
AND3_X1 _13422_ ( .A1(_05962_ ), .A2(\fd_inst[11] ), .A3(_05961_ ), .ZN(_00434_ ) );
AND3_X1 _13423_ ( .A1(_05962_ ), .A2(\fd_inst[10] ), .A3(_05961_ ), .ZN(_00435_ ) );
AND3_X1 _13424_ ( .A1(_05962_ ), .A2(\fd_inst[9] ), .A3(_05961_ ), .ZN(_00436_ ) );
AND3_X1 _13425_ ( .A1(_05962_ ), .A2(\fd_inst[8] ), .A3(_05961_ ), .ZN(_00437_ ) );
AND3_X1 _13426_ ( .A1(_05962_ ), .A2(\fd_inst[7] ), .A3(_05961_ ), .ZN(_00438_ ) );
CLKBUF_X2 _13427_ ( .A(_00637_ ), .Z(_05963_ ) );
AND3_X1 _13428_ ( .A1(_05962_ ), .A2(\fd_inst[6] ), .A3(_05963_ ), .ZN(_00439_ ) );
AND3_X1 _13429_ ( .A1(_05962_ ), .A2(\fd_inst[5] ), .A3(_05963_ ), .ZN(_00440_ ) );
AND3_X1 _13430_ ( .A1(_05962_ ), .A2(\fd_inst[4] ), .A3(_05963_ ), .ZN(_00441_ ) );
AND3_X1 _13431_ ( .A1(_05962_ ), .A2(\fd_inst[3] ), .A3(_05963_ ), .ZN(_00442_ ) );
CLKBUF_X2 _13432_ ( .A(_00863_ ), .Z(_05964_ ) );
AND3_X1 _13433_ ( .A1(_05964_ ), .A2(\fd_inst[2] ), .A3(_05963_ ), .ZN(_00443_ ) );
AND3_X1 _13434_ ( .A1(_05964_ ), .A2(\fd_inst[28] ), .A3(_05963_ ), .ZN(_00444_ ) );
AND3_X1 _13435_ ( .A1(_05964_ ), .A2(\fd_inst[1] ), .A3(_05963_ ), .ZN(_00445_ ) );
AND3_X1 _13436_ ( .A1(_05964_ ), .A2(\fd_inst[0] ), .A3(_05963_ ), .ZN(_00446_ ) );
AND3_X1 _13437_ ( .A1(_05964_ ), .A2(\fd_inst[27] ), .A3(_05963_ ), .ZN(_00447_ ) );
AND3_X1 _13438_ ( .A1(_05964_ ), .A2(\fd_inst[26] ), .A3(_05963_ ), .ZN(_00448_ ) );
CLKBUF_X2 _13439_ ( .A(_00637_ ), .Z(_05965_ ) );
AND3_X1 _13440_ ( .A1(_05964_ ), .A2(\fd_inst[25] ), .A3(_05965_ ), .ZN(_00449_ ) );
AND3_X1 _13441_ ( .A1(_05964_ ), .A2(\fd_inst[24] ), .A3(_05965_ ), .ZN(_00450_ ) );
AND3_X1 _13442_ ( .A1(_05964_ ), .A2(\fd_inst[23] ), .A3(_05965_ ), .ZN(_00451_ ) );
AND3_X1 _13443_ ( .A1(_05964_ ), .A2(\fd_inst[22] ), .A3(_05965_ ), .ZN(_00452_ ) );
NOR4_X1 _13444_ ( .A1(_04463_ ), .A2(fanout_net_3 ), .A3(_04462_ ), .A4(_05391_ ), .ZN(_00453_ ) );
NOR4_X1 _13445_ ( .A1(_04463_ ), .A2(fanout_net_3 ), .A3(_04462_ ), .A4(_05448_ ), .ZN(_00454_ ) );
NOR4_X1 _13446_ ( .A1(_04463_ ), .A2(fanout_net_3 ), .A3(_04462_ ), .A4(_05449_ ), .ZN(_00455_ ) );
BUF_X4 _13447_ ( .A(_00858_ ), .Z(_05966_ ) );
BUF_X4 _13448_ ( .A(_05966_ ), .Z(_05967_ ) );
NOR4_X1 _13449_ ( .A1(_04463_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05450_ ), .ZN(_00456_ ) );
BUF_X4 _13450_ ( .A(_00856_ ), .Z(_05968_ ) );
NOR4_X1 _13451_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05451_ ), .ZN(_00457_ ) );
NOR4_X1 _13452_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05452_ ), .ZN(_00458_ ) );
NOR4_X1 _13453_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05453_ ), .ZN(_00459_ ) );
NOR4_X1 _13454_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05454_ ), .ZN(_00460_ ) );
NOR4_X1 _13455_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05455_ ), .ZN(_00461_ ) );
NOR4_X1 _13456_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05456_ ), .ZN(_00462_ ) );
NOR4_X1 _13457_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05458_ ), .ZN(_00463_ ) );
NOR4_X1 _13458_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05459_ ), .ZN(_00464_ ) );
NOR4_X1 _13459_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05967_ ), .A4(_05460_ ), .ZN(_00465_ ) );
BUF_X4 _13460_ ( .A(_05966_ ), .Z(_05969_ ) );
NOR4_X1 _13461_ ( .A1(_05968_ ), .A2(fanout_net_3 ), .A3(_05969_ ), .A4(_05461_ ), .ZN(_00466_ ) );
BUF_X4 _13462_ ( .A(_00856_ ), .Z(_05970_ ) );
NOR4_X1 _13463_ ( .A1(_05970_ ), .A2(fanout_net_3 ), .A3(_05969_ ), .A4(_05462_ ), .ZN(_00467_ ) );
NOR4_X1 _13464_ ( .A1(_05970_ ), .A2(fanout_net_3 ), .A3(_05969_ ), .A4(_05463_ ), .ZN(_00468_ ) );
NOR4_X1 _13465_ ( .A1(_05970_ ), .A2(fanout_net_3 ), .A3(_05969_ ), .A4(_05464_ ), .ZN(_00469_ ) );
NOR4_X1 _13466_ ( .A1(_05970_ ), .A2(fanout_net_3 ), .A3(_05969_ ), .A4(_05465_ ), .ZN(_00470_ ) );
NOR4_X1 _13467_ ( .A1(_05970_ ), .A2(fanout_net_3 ), .A3(_05969_ ), .A4(_05466_ ), .ZN(_00471_ ) );
NOR4_X1 _13468_ ( .A1(_05970_ ), .A2(fanout_net_4 ), .A3(_05969_ ), .A4(_05467_ ), .ZN(_00472_ ) );
NOR4_X1 _13469_ ( .A1(_05970_ ), .A2(fanout_net_4 ), .A3(_05969_ ), .A4(_05469_ ), .ZN(_00473_ ) );
NOR4_X1 _13470_ ( .A1(_05970_ ), .A2(fanout_net_4 ), .A3(_05969_ ), .A4(_05511_ ), .ZN(_00474_ ) );
NOR4_X1 _13471_ ( .A1(_05970_ ), .A2(fanout_net_4 ), .A3(_05969_ ), .A4(_05496_ ), .ZN(_00475_ ) );
BUF_X4 _13472_ ( .A(_05966_ ), .Z(_05971_ ) );
NOR4_X1 _13473_ ( .A1(_05970_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_05470_ ), .ZN(_00476_ ) );
AND3_X1 _13474_ ( .A1(_05943_ ), .A2(\fc_addr[1] ), .A3(_05965_ ), .ZN(_00477_ ) );
AND3_X1 _13475_ ( .A1(_05943_ ), .A2(\fc_addr[0] ), .A3(_05965_ ), .ZN(_00478_ ) );
BUF_X4 _13476_ ( .A(_00856_ ), .Z(_05972_ ) );
NOR4_X1 _13477_ ( .A1(_05972_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_05471_ ), .ZN(_00479_ ) );
NOR4_X1 _13478_ ( .A1(_05972_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_05472_ ), .ZN(_00480_ ) );
NOR4_X1 _13479_ ( .A1(_05972_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_05473_ ), .ZN(_00481_ ) );
NOR4_X1 _13480_ ( .A1(_05972_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_05474_ ), .ZN(_00482_ ) );
NOR4_X1 _13481_ ( .A1(_05972_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_05475_ ), .ZN(_00483_ ) );
NOR4_X1 _13482_ ( .A1(_05972_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_05476_ ), .ZN(_00484_ ) );
BUF_X4 _13483_ ( .A(_00637_ ), .Z(_05973_ ) );
CLKBUF_X2 _13484_ ( .A(_05973_ ), .Z(_05974_ ) );
AND3_X1 _13485_ ( .A1(_05974_ ), .A2(_00840_ ), .A3(\cf_inst[31] ), .ZN(_00485_ ) );
AND3_X1 _13486_ ( .A1(_05974_ ), .A2(_00840_ ), .A3(\cf_inst[30] ), .ZN(_00486_ ) );
AND3_X1 _13487_ ( .A1(_05974_ ), .A2(_00840_ ), .A3(\cf_inst[21] ), .ZN(_00487_ ) );
AND3_X1 _13488_ ( .A1(_05974_ ), .A2(_00840_ ), .A3(\cf_inst[20] ), .ZN(_00488_ ) );
AND3_X1 _13489_ ( .A1(_05974_ ), .A2(_00840_ ), .A3(\cf_inst[19] ), .ZN(_00489_ ) );
CLKBUF_X2 _13490_ ( .A(_00772_ ), .Z(_05975_ ) );
AND3_X1 _13491_ ( .A1(_05974_ ), .A2(_05975_ ), .A3(\cf_inst[18] ), .ZN(_00490_ ) );
AND3_X1 _13492_ ( .A1(_05974_ ), .A2(_05975_ ), .A3(\cf_inst[17] ), .ZN(_00491_ ) );
AND3_X1 _13493_ ( .A1(_05974_ ), .A2(_05975_ ), .A3(\cf_inst[16] ), .ZN(_00492_ ) );
AND3_X1 _13494_ ( .A1(_05974_ ), .A2(_05975_ ), .A3(\cf_inst[15] ), .ZN(_00493_ ) );
AND3_X1 _13495_ ( .A1(_05974_ ), .A2(_05975_ ), .A3(\cf_inst[14] ), .ZN(_00494_ ) );
CLKBUF_X2 _13496_ ( .A(_05973_ ), .Z(_05976_ ) );
AND3_X1 _13497_ ( .A1(_05976_ ), .A2(_05975_ ), .A3(\cf_inst[13] ), .ZN(_00495_ ) );
AND3_X1 _13498_ ( .A1(_05976_ ), .A2(_05975_ ), .A3(\cf_inst[12] ), .ZN(_00496_ ) );
AND3_X1 _13499_ ( .A1(_05976_ ), .A2(_05975_ ), .A3(\cf_inst[29] ), .ZN(_00497_ ) );
AND3_X1 _13500_ ( .A1(_05976_ ), .A2(_05975_ ), .A3(\cf_inst[11] ), .ZN(_00498_ ) );
AND3_X1 _13501_ ( .A1(_05976_ ), .A2(_05975_ ), .A3(\cf_inst[10] ), .ZN(_00499_ ) );
CLKBUF_X2 _13502_ ( .A(_00772_ ), .Z(_05977_ ) );
AND3_X1 _13503_ ( .A1(_05976_ ), .A2(_05977_ ), .A3(\cf_inst[9] ), .ZN(_00500_ ) );
AND3_X1 _13504_ ( .A1(_05976_ ), .A2(_05977_ ), .A3(\cf_inst[8] ), .ZN(_00501_ ) );
AND3_X1 _13505_ ( .A1(_05976_ ), .A2(_05977_ ), .A3(\cf_inst[7] ), .ZN(_00502_ ) );
AND3_X1 _13506_ ( .A1(_05976_ ), .A2(_05977_ ), .A3(\cf_inst[6] ), .ZN(_00503_ ) );
AND3_X1 _13507_ ( .A1(_05976_ ), .A2(_05977_ ), .A3(\cf_inst[5] ), .ZN(_00504_ ) );
CLKBUF_X2 _13508_ ( .A(_05973_ ), .Z(_05978_ ) );
AND3_X1 _13509_ ( .A1(_05978_ ), .A2(_05977_ ), .A3(\cf_inst[4] ), .ZN(_00505_ ) );
AND3_X1 _13510_ ( .A1(_05978_ ), .A2(_05977_ ), .A3(\cf_inst[3] ), .ZN(_00506_ ) );
AND3_X1 _13511_ ( .A1(_05978_ ), .A2(_05977_ ), .A3(\cf_inst[2] ), .ZN(_00507_ ) );
AND3_X1 _13512_ ( .A1(_05978_ ), .A2(_05977_ ), .A3(\cf_inst[28] ), .ZN(_00508_ ) );
AND3_X1 _13513_ ( .A1(_05978_ ), .A2(_05977_ ), .A3(\cf_inst[1] ), .ZN(_00509_ ) );
AND3_X1 _13514_ ( .A1(_05978_ ), .A2(_00779_ ), .A3(\cf_inst[0] ), .ZN(_00510_ ) );
AND3_X1 _13515_ ( .A1(_05978_ ), .A2(_00779_ ), .A3(\cf_inst[27] ), .ZN(_00511_ ) );
AND3_X1 _13516_ ( .A1(_05978_ ), .A2(_00779_ ), .A3(\cf_inst[26] ), .ZN(_00512_ ) );
AND3_X1 _13517_ ( .A1(_05978_ ), .A2(_00779_ ), .A3(\cf_inst[25] ), .ZN(_00513_ ) );
AND3_X1 _13518_ ( .A1(_05978_ ), .A2(_00779_ ), .A3(\cf_inst[24] ), .ZN(_00514_ ) );
AND3_X1 _13519_ ( .A1(_00866_ ), .A2(_00779_ ), .A3(\cf_inst[23] ), .ZN(_00515_ ) );
AND3_X1 _13520_ ( .A1(_00866_ ), .A2(_00779_ ), .A3(\cf_inst[22] ), .ZN(_00516_ ) );
NAND2_X1 _13521_ ( .A1(_05836_ ), .A2(_05837_ ), .ZN(_05979_ ) );
NOR2_X1 _13522_ ( .A1(_05979_ ), .A2(_05952_ ), .ZN(\u_icache.cready_$_ANDNOT__A_Y ) );
AND4_X1 _13523_ ( .A1(ifu_ready ), .A2(_05836_ ), .A3(_00873_ ), .A4(_05837_ ), .ZN(_00517_ ) );
AOI211_X1 _13524_ ( .A(_00767_ ), .B(_04456_ ), .C1(_00760_ ), .C2(_00761_ ), .ZN(_00518_ ) );
AND3_X1 _13525_ ( .A1(_01536_ ), .A2(_05966_ ), .A3(_01552_ ), .ZN(_05980_ ) );
AOI211_X1 _13526_ ( .A(_00771_ ), .B(_04585_ ), .C1(_04588_ ), .C2(_04645_ ), .ZN(_05981_ ) );
AND3_X4 _13527_ ( .A1(\fc_addr[4] ), .A2(\fc_addr[3] ), .A3(\fc_addr[2] ), .ZN(_05982_ ) );
AND2_X1 _13528_ ( .A1(_05982_ ), .A2(\fc_addr[5] ), .ZN(_05983_ ) );
AND2_X2 _13529_ ( .A1(_05983_ ), .A2(\fc_addr[6] ), .ZN(_05984_ ) );
AND2_X1 _13530_ ( .A1(_05984_ ), .A2(\fc_addr[7] ), .ZN(_05985_ ) );
AND2_X1 _13531_ ( .A1(_05985_ ), .A2(\fc_addr[8] ), .ZN(_05986_ ) );
AND2_X4 _13532_ ( .A1(_05986_ ), .A2(\fc_addr[9] ), .ZN(_05987_ ) );
AND2_X1 _13533_ ( .A1(_05987_ ), .A2(\fc_addr[10] ), .ZN(_05988_ ) );
AND2_X1 _13534_ ( .A1(_05988_ ), .A2(\fc_addr[11] ), .ZN(_05989_ ) );
AND2_X1 _13535_ ( .A1(_05989_ ), .A2(\fc_addr[12] ), .ZN(_05990_ ) );
AND2_X1 _13536_ ( .A1(_05990_ ), .A2(\fc_addr[13] ), .ZN(_05991_ ) );
AND2_X1 _13537_ ( .A1(_05991_ ), .A2(\fc_addr[14] ), .ZN(_05992_ ) );
AND2_X1 _13538_ ( .A1(_05992_ ), .A2(\fc_addr[15] ), .ZN(_05993_ ) );
AND2_X1 _13539_ ( .A1(_05993_ ), .A2(\fc_addr[16] ), .ZN(_05994_ ) );
AND2_X1 _13540_ ( .A1(_05994_ ), .A2(\fc_addr[17] ), .ZN(_05995_ ) );
AND2_X1 _13541_ ( .A1(_05995_ ), .A2(\fc_addr[18] ), .ZN(_05996_ ) );
AND2_X1 _13542_ ( .A1(_05996_ ), .A2(\fc_addr[19] ), .ZN(_05997_ ) );
AND3_X1 _13543_ ( .A1(_05997_ ), .A2(\fc_addr[21] ), .A3(\fc_addr[20] ), .ZN(_05998_ ) );
AND3_X4 _13544_ ( .A1(_05998_ ), .A2(\fc_addr[23] ), .A3(\fc_addr[22] ), .ZN(_05999_ ) );
AND2_X1 _13545_ ( .A1(_05999_ ), .A2(\fc_addr[24] ), .ZN(_06000_ ) );
AND2_X1 _13546_ ( .A1(_06000_ ), .A2(\fc_addr[25] ), .ZN(_06001_ ) );
AND3_X4 _13547_ ( .A1(_06001_ ), .A2(\fc_addr[27] ), .A3(\fc_addr[26] ), .ZN(_06002_ ) );
AND3_X1 _13548_ ( .A1(_06002_ ), .A2(\fc_addr[29] ), .A3(\fc_addr[28] ), .ZN(_06003_ ) );
XNOR2_X1 _13549_ ( .A(_06003_ ), .B(_05448_ ), .ZN(_06004_ ) );
AOI21_X1 _13550_ ( .A(_05981_ ), .B1(_06004_ ), .B2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06005_ ) );
BUF_X4 _13551_ ( .A(_05973_ ), .Z(_06006_ ) );
AOI211_X1 _13552_ ( .A(fanout_net_4 ), .B(_05980_ ), .C1(_06005_ ), .C2(_06006_ ), .ZN(_00519_ ) );
AND3_X1 _13553_ ( .A1(_02209_ ), .A2(_05966_ ), .A3(_02215_ ), .ZN(_06007_ ) );
BUF_X4 _13554_ ( .A(_00770_ ), .Z(_06008_ ) );
BUF_X4 _13555_ ( .A(_06008_ ), .Z(_06009_ ) );
AOI21_X1 _13556_ ( .A(\fc_addr[29] ), .B1(_06002_ ), .B2(\fc_addr[28] ), .ZN(_06010_ ) );
OAI21_X1 _13557_ ( .A(_06009_ ), .B1(_06003_ ), .B2(_06010_ ), .ZN(_06011_ ) );
OAI21_X1 _13558_ ( .A(_06011_ ), .B1(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .B2(_05011_ ), .ZN(_06012_ ) );
AOI211_X1 _13559_ ( .A(fanout_net_4 ), .B(_06007_ ), .C1(_06012_ ), .C2(_06006_ ), .ZN(_00520_ ) );
AND3_X1 _13560_ ( .A1(_01696_ ), .A2(_05966_ ), .A3(_01714_ ), .ZN(_06013_ ) );
INV_X1 _13561_ ( .A(_05997_ ), .ZN(_06014_ ) );
OAI21_X1 _13562_ ( .A(_06008_ ), .B1(_06014_ ), .B2(_05450_ ), .ZN(_06015_ ) );
AOI21_X1 _13563_ ( .A(_06015_ ), .B1(_05450_ ), .B2(_06014_ ), .ZN(_06016_ ) );
AOI21_X1 _13564_ ( .A(_06016_ ), .B1(_04756_ ), .B2(_05959_ ), .ZN(_06017_ ) );
AOI211_X1 _13565_ ( .A(fanout_net_4 ), .B(_06013_ ), .C1(_06017_ ), .C2(_06006_ ), .ZN(_00521_ ) );
BUF_X4 _13566_ ( .A(_00858_ ), .Z(_06018_ ) );
AOI211_X1 _13567_ ( .A(_06008_ ), .B(_04757_ ), .C1(_04765_ ), .C2(_04796_ ), .ZN(_06019_ ) );
NAND4_X1 _13568_ ( .A1(\fc_addr[17] ), .A2(\fc_addr[16] ), .A3(\fc_addr[15] ), .A4(\fc_addr[14] ), .ZN(_06020_ ) );
NAND2_X1 _13569_ ( .A1(\fc_addr[11] ), .A2(\fc_addr[10] ), .ZN(_06021_ ) );
NOR4_X1 _13570_ ( .A1(_06020_ ), .A2(_06021_ ), .A3(_05458_ ), .A4(_05459_ ), .ZN(_06022_ ) );
NAND3_X1 _13571_ ( .A1(_05987_ ), .A2(\fc_addr[18] ), .A3(_06022_ ), .ZN(_06023_ ) );
XNOR2_X1 _13572_ ( .A(_06023_ ), .B(\fc_addr[19] ), .ZN(_06024_ ) );
AOI211_X1 _13573_ ( .A(_06018_ ), .B(_06019_ ), .C1(_06009_ ), .C2(_06024_ ), .ZN(_06025_ ) );
BUF_X4 _13574_ ( .A(_00859_ ), .Z(_06026_ ) );
AOI211_X1 _13575_ ( .A(fanout_net_4 ), .B(_06025_ ), .C1(_06026_ ), .C2(_01790_ ), .ZN(_00522_ ) );
AOI211_X1 _13576_ ( .A(_06008_ ), .B(_04797_ ), .C1(_04799_ ), .C2(_04833_ ), .ZN(_06027_ ) );
NAND2_X1 _13577_ ( .A1(_05987_ ), .A2(_06022_ ), .ZN(_06028_ ) );
XNOR2_X1 _13578_ ( .A(_06028_ ), .B(\fc_addr[18] ), .ZN(_06029_ ) );
AOI211_X1 _13579_ ( .A(_06018_ ), .B(_06027_ ), .C1(_06009_ ), .C2(_06029_ ), .ZN(_06030_ ) );
AOI211_X1 _13580_ ( .A(fanout_net_4 ), .B(_06030_ ), .C1(_06026_ ), .C2(_01879_ ), .ZN(_00523_ ) );
AOI211_X1 _13581_ ( .A(_06008_ ), .B(_04834_ ), .C1(_04837_ ), .C2(_04866_ ), .ZN(_06031_ ) );
XNOR2_X1 _13582_ ( .A(_05994_ ), .B(_05453_ ), .ZN(_06032_ ) );
AOI211_X1 _13583_ ( .A(_06018_ ), .B(_06031_ ), .C1(_06009_ ), .C2(_06032_ ), .ZN(_06033_ ) );
AOI211_X1 _13584_ ( .A(fanout_net_4 ), .B(_06033_ ), .C1(_06026_ ), .C2(_01934_ ), .ZN(_00524_ ) );
AOI211_X1 _13585_ ( .A(_06008_ ), .B(_04867_ ), .C1(_04883_ ), .C2(_04886_ ), .ZN(_06034_ ) );
XNOR2_X1 _13586_ ( .A(_05993_ ), .B(_05454_ ), .ZN(_06035_ ) );
AOI211_X1 _13587_ ( .A(_06018_ ), .B(_06034_ ), .C1(_06009_ ), .C2(_06035_ ), .ZN(_06036_ ) );
AOI211_X1 _13588_ ( .A(fanout_net_4 ), .B(_06036_ ), .C1(_06026_ ), .C2(_01990_ ), .ZN(_00525_ ) );
INV_X1 _13589_ ( .A(_05992_ ), .ZN(_06037_ ) );
OAI21_X1 _13590_ ( .A(_06008_ ), .B1(_06037_ ), .B2(_05455_ ), .ZN(_06038_ ) );
AOI21_X1 _13591_ ( .A(_06038_ ), .B1(_05455_ ), .B2(_06037_ ), .ZN(_06039_ ) );
AOI21_X1 _13592_ ( .A(_04887_ ), .B1(_04897_ ), .B2(_04918_ ), .ZN(_06040_ ) );
AOI211_X1 _13593_ ( .A(_06018_ ), .B(_06039_ ), .C1(_06040_ ), .C2(_05959_ ), .ZN(_06041_ ) );
AOI211_X1 _13594_ ( .A(fanout_net_4 ), .B(_06041_ ), .C1(_06026_ ), .C2(_02031_ ), .ZN(_00526_ ) );
INV_X1 _13595_ ( .A(_05991_ ), .ZN(_06042_ ) );
OAI21_X1 _13596_ ( .A(_00770_ ), .B1(_06042_ ), .B2(_05456_ ), .ZN(_06043_ ) );
AOI21_X1 _13597_ ( .A(_06043_ ), .B1(_05456_ ), .B2(_06042_ ), .ZN(_06044_ ) );
AOI21_X1 _13598_ ( .A(_04919_ ), .B1(_04921_ ), .B2(_04940_ ), .ZN(_06045_ ) );
BUF_X4 _13599_ ( .A(_05958_ ), .Z(_06046_ ) );
AOI211_X1 _13600_ ( .A(_06018_ ), .B(_06044_ ), .C1(_06045_ ), .C2(_06046_ ), .ZN(_06047_ ) );
AOI211_X1 _13601_ ( .A(fanout_net_4 ), .B(_06047_ ), .C1(_06026_ ), .C2(_02085_ ), .ZN(_00527_ ) );
INV_X1 _13602_ ( .A(_05990_ ), .ZN(_06048_ ) );
OAI21_X1 _13603_ ( .A(_00770_ ), .B1(_06048_ ), .B2(_05458_ ), .ZN(_06049_ ) );
AOI21_X1 _13604_ ( .A(_06049_ ), .B1(_05458_ ), .B2(_06048_ ), .ZN(_06050_ ) );
AOI21_X1 _13605_ ( .A(_04941_ ), .B1(_04944_ ), .B2(_04967_ ), .ZN(_06051_ ) );
AOI211_X1 _13606_ ( .A(_06018_ ), .B(_06050_ ), .C1(_06051_ ), .C2(_06046_ ), .ZN(_06052_ ) );
AOI211_X1 _13607_ ( .A(fanout_net_4 ), .B(_06052_ ), .C1(_06026_ ), .C2(_02131_ ), .ZN(_00528_ ) );
INV_X1 _13608_ ( .A(_05989_ ), .ZN(_06053_ ) );
OAI21_X1 _13609_ ( .A(_00770_ ), .B1(_06053_ ), .B2(_05459_ ), .ZN(_06054_ ) );
AOI21_X1 _13610_ ( .A(_06054_ ), .B1(_05459_ ), .B2(_06053_ ), .ZN(_06055_ ) );
AOI211_X1 _13611_ ( .A(_06018_ ), .B(_06055_ ), .C1(_04988_ ), .C2(_06046_ ), .ZN(_06056_ ) );
AOI211_X1 _13612_ ( .A(fanout_net_4 ), .B(_06056_ ), .C1(_06026_ ), .C2(_02182_ ), .ZN(_00529_ ) );
AND3_X1 _13613_ ( .A1(_02256_ ), .A2(_05966_ ), .A3(_02262_ ), .ZN(_06057_ ) );
INV_X1 _13614_ ( .A(_05988_ ), .ZN(_06058_ ) );
OAI21_X1 _13615_ ( .A(_06008_ ), .B1(_06058_ ), .B2(_05461_ ), .ZN(_06059_ ) );
AOI21_X1 _13616_ ( .A(_06059_ ), .B1(_05461_ ), .B2(_06058_ ), .ZN(_06060_ ) );
AOI21_X1 _13617_ ( .A(_05012_ ), .B1(_05021_ ), .B2(_05042_ ), .ZN(_06061_ ) );
AOI21_X1 _13618_ ( .A(_06060_ ), .B1(_06061_ ), .B2(_05959_ ), .ZN(_06062_ ) );
AOI211_X1 _13619_ ( .A(fanout_net_4 ), .B(_06057_ ), .C1(_06062_ ), .C2(_06006_ ), .ZN(_00530_ ) );
AND3_X1 _13620_ ( .A1(_02722_ ), .A2(_05966_ ), .A3(_02728_ ), .ZN(_06063_ ) );
AOI211_X1 _13621_ ( .A(_00771_ ), .B(_05234_ ), .C1(_05236_ ), .C2(_05254_ ), .ZN(_06064_ ) );
XNOR2_X1 _13622_ ( .A(_06002_ ), .B(_05470_ ), .ZN(_06065_ ) );
AOI21_X1 _13623_ ( .A(_06064_ ), .B1(_06065_ ), .B2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06066_ ) );
AOI211_X1 _13624_ ( .A(fanout_net_4 ), .B(_06063_ ), .C1(_06066_ ), .C2(_06006_ ), .ZN(_00531_ ) );
INV_X1 _13625_ ( .A(_05987_ ), .ZN(_06067_ ) );
OAI21_X1 _13626_ ( .A(_00770_ ), .B1(_06067_ ), .B2(_05462_ ), .ZN(_06068_ ) );
AOI21_X1 _13627_ ( .A(_06068_ ), .B1(_05462_ ), .B2(_06067_ ), .ZN(_06069_ ) );
AOI21_X1 _13628_ ( .A(_05043_ ), .B1(_05045_ ), .B2(_05066_ ), .ZN(_06070_ ) );
AOI211_X1 _13629_ ( .A(_06018_ ), .B(_06069_ ), .C1(_06070_ ), .C2(_06046_ ), .ZN(_06071_ ) );
AOI211_X1 _13630_ ( .A(fanout_net_4 ), .B(_06071_ ), .C1(_06026_ ), .C2(_02310_ ), .ZN(_00532_ ) );
AND3_X1 _13631_ ( .A1(_02350_ ), .A2(_05966_ ), .A3(_02355_ ), .ZN(_06072_ ) );
INV_X1 _13632_ ( .A(_05986_ ), .ZN(_06073_ ) );
OAI21_X1 _13633_ ( .A(_06008_ ), .B1(_06073_ ), .B2(_05463_ ), .ZN(_06074_ ) );
AOI21_X1 _13634_ ( .A(_06074_ ), .B1(_05463_ ), .B2(_06073_ ), .ZN(_06075_ ) );
AOI21_X1 _13635_ ( .A(_05067_ ), .B1(_05070_ ), .B2(_05090_ ), .ZN(_06076_ ) );
AOI21_X1 _13636_ ( .A(_06075_ ), .B1(_06076_ ), .B2(_05959_ ), .ZN(_06077_ ) );
AOI211_X1 _13637_ ( .A(fanout_net_4 ), .B(_06072_ ), .C1(_06077_ ), .C2(_06006_ ), .ZN(_00533_ ) );
AND3_X1 _13638_ ( .A1(_02395_ ), .A2(_05966_ ), .A3(_02401_ ), .ZN(_06078_ ) );
XNOR2_X1 _13639_ ( .A(_05985_ ), .B(\fc_addr[8] ), .ZN(_06079_ ) );
MUX2_X1 _13640_ ( .A(_06079_ ), .B(_05110_ ), .S(_06046_ ), .Z(_06080_ ) );
AOI211_X1 _13641_ ( .A(fanout_net_4 ), .B(_06078_ ), .C1(_06080_ ), .C2(_06006_ ), .ZN(_00534_ ) );
AND3_X1 _13642_ ( .A1(_04057_ ), .A2(_06018_ ), .A3(_04058_ ), .ZN(_06081_ ) );
XNOR2_X1 _13643_ ( .A(_05984_ ), .B(\fc_addr[7] ), .ZN(_06082_ ) );
MUX2_X1 _13644_ ( .A(_06082_ ), .B(_05137_ ), .S(_06046_ ), .Z(_06083_ ) );
AOI211_X1 _13645_ ( .A(fanout_net_4 ), .B(_06081_ ), .C1(_06006_ ), .C2(_06083_ ), .ZN(_00535_ ) );
NAND2_X1 _13646_ ( .A1(_00858_ ), .A2(_00772_ ), .ZN(_06084_ ) );
BUF_X4 _13647_ ( .A(_06084_ ), .Z(_06085_ ) );
AOI21_X1 _13648_ ( .A(\fc_addr[6] ), .B1(_05982_ ), .B2(\fc_addr[5] ), .ZN(_06086_ ) );
NOR3_X1 _13649_ ( .A1(_05984_ ), .A2(_06046_ ), .A3(_06086_ ), .ZN(_06087_ ) );
AOI21_X1 _13650_ ( .A(_06087_ ), .B1(_05157_ ), .B2(_05959_ ), .ZN(_06088_ ) );
OAI22_X1 _13651_ ( .A1(_02485_ ), .A2(_06085_ ), .B1(_04456_ ), .B2(_06088_ ), .ZN(_00536_ ) );
INV_X1 _13652_ ( .A(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B ), .ZN(_06089_ ) );
AOI21_X1 _13653_ ( .A(\fc_addr[5] ), .B1(_05502_ ), .B2(_06089_ ), .ZN(_06090_ ) );
AND4_X1 _13654_ ( .A1(\fc_addr[5] ), .A2(_06089_ ), .A3(\fc_addr[3] ), .A4(\fc_addr[2] ), .ZN(_06091_ ) );
NOR3_X1 _13655_ ( .A1(_06090_ ), .A2(_06091_ ), .A3(_06046_ ), .ZN(_06092_ ) );
AOI21_X1 _13656_ ( .A(_06092_ ), .B1(_05178_ ), .B2(_05959_ ), .ZN(_06093_ ) );
OAI22_X1 _13657_ ( .A1(_02527_ ), .A2(_06085_ ), .B1(_04456_ ), .B2(_06093_ ), .ZN(_00537_ ) );
AOI21_X1 _13658_ ( .A(\fc_addr[4] ), .B1(\fc_addr[3] ), .B2(\fc_addr[2] ), .ZN(_06094_ ) );
NOR3_X1 _13659_ ( .A1(_05958_ ), .A2(_05982_ ), .A3(_06094_ ), .ZN(_06095_ ) );
AOI21_X1 _13660_ ( .A(_05179_ ), .B1(_05193_ ), .B2(_05195_ ), .ZN(_06096_ ) );
AOI21_X1 _13661_ ( .A(_06095_ ), .B1(_06096_ ), .B2(_06046_ ), .ZN(_06097_ ) );
MUX2_X1 _13662_ ( .A(_06097_ ), .B(_02573_ ), .S(_00858_ ), .Z(_06098_ ) );
NOR2_X1 _13663_ ( .A1(_06098_ ), .A2(fanout_net_4 ), .ZN(_00538_ ) );
XNOR2_X1 _13664_ ( .A(\fc_addr[3] ), .B(\fc_addr[2] ), .ZN(_06099_ ) );
MUX2_X1 _13665_ ( .A(_06099_ ), .B(_05216_ ), .S(_06046_ ), .Z(_06100_ ) );
OAI22_X1 _13666_ ( .A1(_02631_ ), .A2(_06085_ ), .B1(_04456_ ), .B2(_06100_ ), .ZN(_00539_ ) );
OAI21_X1 _13667_ ( .A(_00779_ ), .B1(_00000_ ), .B2(\fc_addr[4] ), .ZN(_06101_ ) );
AOI21_X1 _13668_ ( .A(_06101_ ), .B1(_06098_ ), .B2(_00000_ ), .ZN(_00540_ ) );
AOI211_X1 _13669_ ( .A(_00771_ ), .B(_05217_ ), .C1(_05231_ ), .C2(_05233_ ), .ZN(_06102_ ) );
AOI21_X1 _13670_ ( .A(_06102_ ), .B1(\u_ifu.pc_$_SDFFE_PP0N__Q_28_D_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06009_ ), .ZN(_06103_ ) );
OAI22_X1 _13671_ ( .A1(_02684_ ), .A2(_06085_ ), .B1(_06103_ ), .B2(_04456_ ), .ZN(_00541_ ) );
AOI21_X1 _13672_ ( .A(\fc_addr[27] ), .B1(_06001_ ), .B2(\fc_addr[26] ), .ZN(_06104_ ) );
OAI21_X1 _13673_ ( .A(_00771_ ), .B1(_06002_ ), .B2(_06104_ ), .ZN(_06105_ ) );
OAI211_X1 _13674_ ( .A(_00873_ ), .B(_06105_ ), .C1(_05298_ ), .C2(_06009_ ), .ZN(_06106_ ) );
AND2_X1 _13675_ ( .A1(_02858_ ), .A2(_02864_ ), .ZN(_06107_ ) );
OAI21_X1 _13676_ ( .A(_06106_ ), .B1(_06107_ ), .B2(_06085_ ), .ZN(_00542_ ) );
AND2_X1 _13677_ ( .A1(_06001_ ), .A2(\fc_addr[26] ), .ZN(_06108_ ) );
AOI21_X1 _13678_ ( .A(\fc_addr[26] ), .B1(_06000_ ), .B2(\fc_addr[25] ), .ZN(_06109_ ) );
OAI21_X1 _13679_ ( .A(_06009_ ), .B1(_06108_ ), .B2(_06109_ ), .ZN(_06110_ ) );
OAI211_X1 _13680_ ( .A(_06110_ ), .B(_00873_ ), .C1(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .C2(_05315_ ), .ZN(_06111_ ) );
AND2_X1 _13681_ ( .A1(_02897_ ), .A2(_02902_ ), .ZN(_06112_ ) );
OAI21_X1 _13682_ ( .A(_06111_ ), .B1(_06112_ ), .B2(_06085_ ), .ZN(_00543_ ) );
AOI21_X1 _13683_ ( .A(\fc_addr[25] ), .B1(_05999_ ), .B2(\fc_addr[24] ), .ZN(_06113_ ) );
OAI21_X1 _13684_ ( .A(_00771_ ), .B1(_06001_ ), .B2(_06113_ ), .ZN(_06114_ ) );
OAI211_X1 _13685_ ( .A(_00873_ ), .B(_06114_ ), .C1(_05337_ ), .C2(_06009_ ), .ZN(_06115_ ) );
AND2_X1 _13686_ ( .A1(_02935_ ), .A2(_02940_ ), .ZN(_06116_ ) );
OAI21_X1 _13687_ ( .A(_06115_ ), .B1(_06116_ ), .B2(_06085_ ), .ZN(_00544_ ) );
INV_X1 _13688_ ( .A(_05999_ ), .ZN(_06117_ ) );
OAI21_X1 _13689_ ( .A(_06008_ ), .B1(_06117_ ), .B2(_05474_ ), .ZN(_06118_ ) );
AOI21_X1 _13690_ ( .A(_06118_ ), .B1(_05474_ ), .B2(_06117_ ), .ZN(_06119_ ) );
AOI21_X1 _13691_ ( .A(_06119_ ), .B1(_05959_ ), .B2(_05354_ ), .ZN(_06120_ ) );
BUF_X4 _13692_ ( .A(_00874_ ), .Z(_06121_ ) );
OAI22_X1 _13693_ ( .A1(_06120_ ), .A2(_06121_ ), .B1(_02979_ ), .B2(_06085_ ), .ZN(_00545_ ) );
AOI211_X1 _13694_ ( .A(_00771_ ), .B(_05355_ ), .C1(_05361_ ), .C2(_05373_ ), .ZN(_06122_ ) );
AND2_X1 _13695_ ( .A1(_05998_ ), .A2(\fc_addr[22] ), .ZN(_06123_ ) );
XNOR2_X1 _13696_ ( .A(_06123_ ), .B(_05475_ ), .ZN(_06124_ ) );
AOI21_X1 _13697_ ( .A(_06122_ ), .B1(_06124_ ), .B2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06125_ ) );
AND2_X1 _13698_ ( .A1(_03013_ ), .A2(_03018_ ), .ZN(_06126_ ) );
OAI22_X1 _13699_ ( .A1(_06125_ ), .A2(_06121_ ), .B1(_06126_ ), .B2(_06085_ ), .ZN(_00546_ ) );
AOI211_X1 _13700_ ( .A(_00771_ ), .B(_05374_ ), .C1(_05376_ ), .C2(_05389_ ), .ZN(_06127_ ) );
XNOR2_X1 _13701_ ( .A(_05998_ ), .B(_05476_ ), .ZN(_06128_ ) );
AOI21_X1 _13702_ ( .A(_06127_ ), .B1(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .B2(_06128_ ), .ZN(_06129_ ) );
OAI22_X1 _13703_ ( .A1(_06129_ ), .A2(_06121_ ), .B1(_03063_ ), .B2(_06084_ ), .ZN(_00547_ ) );
AOI211_X1 _13704_ ( .A(_00771_ ), .B(_04646_ ), .C1(_04653_ ), .C2(_04711_ ), .ZN(_06130_ ) );
NOR3_X1 _13705_ ( .A1(_06028_ ), .A2(_05451_ ), .A3(_05452_ ), .ZN(_06131_ ) );
NAND2_X1 _13706_ ( .A1(_06131_ ), .A2(\fc_addr[20] ), .ZN(_06132_ ) );
XNOR2_X1 _13707_ ( .A(_06132_ ), .B(\fc_addr[21] ), .ZN(_06133_ ) );
AOI21_X1 _13708_ ( .A(_06130_ ), .B1(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .B2(_06133_ ), .ZN(_06134_ ) );
OAI22_X1 _13709_ ( .A1(_06134_ ), .A2(_06121_ ), .B1(_01635_ ), .B2(_06084_ ), .ZN(_00548_ ) );
NAND3_X1 _13710_ ( .A1(_00637_ ), .A2(_00772_ ), .A3(_05958_ ), .ZN(_06135_ ) );
OR3_X1 _13711_ ( .A1(_05272_ ), .A2(_05273_ ), .A3(_06135_ ), .ZN(_06136_ ) );
OAI21_X1 _13712_ ( .A(_06136_ ), .B1(_02769_ ), .B2(_06085_ ), .ZN(_00549_ ) );
OAI22_X1 _13713_ ( .A1(_04219_ ), .A2(_06135_ ), .B1(_02817_ ), .B2(_06084_ ), .ZN(_00550_ ) );
AND2_X1 _13714_ ( .A1(_01422_ ), .A2(_01445_ ), .ZN(_06137_ ) );
OAI21_X1 _13715_ ( .A(_05973_ ), .B1(_04579_ ), .B2(_06009_ ), .ZN(_06138_ ) );
AND3_X1 _13716_ ( .A1(_06003_ ), .A2(_05391_ ), .A3(\fc_addr[30] ), .ZN(_06139_ ) );
AOI21_X1 _13717_ ( .A(_05391_ ), .B1(_06003_ ), .B2(\fc_addr[30] ), .ZN(_06140_ ) );
NOR3_X1 _13718_ ( .A1(_06139_ ), .A2(_06140_ ), .A3(_05959_ ), .ZN(_06141_ ) );
OAI221_X1 _13719_ ( .A(_00774_ ), .B1(_06006_ ), .B2(_06137_ ), .C1(_06138_ ), .C2(_06141_ ), .ZN(_00551_ ) );
OR2_X1 _13720_ ( .A1(_01217_ ), .A2(\u_lsu.reading ), .ZN(_06142_ ) );
NOR4_X1 _13721_ ( .A1(_05972_ ), .A2(fanout_net_4 ), .A3(_05971_ ), .A4(_06142_ ), .ZN(_00552_ ) );
OAI21_X1 _13722_ ( .A(\u_arbiter.wvalid ), .B1(_01143_ ), .B2(\u_arbiter.working ), .ZN(_06143_ ) );
NOR4_X1 _13723_ ( .A1(_06121_ ), .A2(\u_lsu.writing ), .A3(_00879_ ), .A4(_06143_ ), .ZN(_00553_ ) );
AND2_X1 _13724_ ( .A1(\u_lsu.rcount[1] ), .A2(\u_lsu.rcount[0] ), .ZN(_06144_ ) );
AND2_X1 _13725_ ( .A1(_06144_ ), .A2(\u_lsu.rcount[2] ), .ZN(_06145_ ) );
AND2_X1 _13726_ ( .A1(_06145_ ), .A2(\u_lsu.rcount[3] ), .ZN(_06146_ ) );
AND2_X1 _13727_ ( .A1(_06146_ ), .A2(\u_lsu.rcount[4] ), .ZN(_06147_ ) );
AND2_X1 _13728_ ( .A1(_06147_ ), .A2(\u_lsu.rcount[5] ), .ZN(_06148_ ) );
AND2_X1 _13729_ ( .A1(_06148_ ), .A2(\u_lsu.rcount[6] ), .ZN(_06149_ ) );
XNOR2_X1 _13730_ ( .A(_06149_ ), .B(\u_lsu.rcount[7] ), .ZN(_06150_ ) );
NOR3_X1 _13731_ ( .A1(_06150_ ), .A2(_04455_ ), .A3(_04456_ ), .ZN(_00554_ ) );
OAI211_X1 _13732_ ( .A(_05965_ ), .B(_05943_ ), .C1(\u_lsu.rcount[6] ), .C2(_06148_ ), .ZN(_06151_ ) );
NOR2_X1 _13733_ ( .A1(_06151_ ), .A2(_06149_ ), .ZN(_00555_ ) );
OAI211_X1 _13734_ ( .A(_05965_ ), .B(_05943_ ), .C1(\u_lsu.rcount[5] ), .C2(_06147_ ), .ZN(_06152_ ) );
NOR2_X1 _13735_ ( .A1(_06152_ ), .A2(_06148_ ), .ZN(_00556_ ) );
OAI211_X1 _13736_ ( .A(_05965_ ), .B(_00864_ ), .C1(\u_lsu.rcount[4] ), .C2(_06146_ ), .ZN(_06153_ ) );
NOR2_X1 _13737_ ( .A1(_06153_ ), .A2(_06147_ ), .ZN(_00557_ ) );
OAI211_X1 _13738_ ( .A(_05973_ ), .B(_00864_ ), .C1(\u_lsu.rcount[3] ), .C2(_06145_ ), .ZN(_06154_ ) );
NOR2_X1 _13739_ ( .A1(_06154_ ), .A2(_06146_ ), .ZN(_00558_ ) );
NOR2_X1 _13740_ ( .A1(\u_lsu.rcount[1] ), .A2(\u_lsu.rcount[0] ), .ZN(_06155_ ) );
MUX2_X1 _13741_ ( .A(_06155_ ), .B(_06144_ ), .S(_01195_ ), .Z(_06156_ ) );
OR4_X1 _13742_ ( .A1(\u_lsu.rcount[4] ), .A2(\u_lsu.rcount[3] ), .A3(\u_lsu.rcount[2] ), .A4(\u_lsu.rcount[7] ), .ZN(_06157_ ) );
NOR3_X1 _13743_ ( .A1(_06157_ ), .A2(\u_lsu.rcount[6] ), .A3(\u_lsu.rcount[5] ), .ZN(_06158_ ) );
AND2_X1 _13744_ ( .A1(_06156_ ), .A2(_06158_ ), .ZN(_06159_ ) );
AOI21_X1 _13745_ ( .A(\u_lsu.rcount[2] ), .B1(\u_lsu.rcount[1] ), .B2(\u_lsu.rcount[0] ), .ZN(_06160_ ) );
NOR4_X1 _13746_ ( .A1(_04467_ ), .A2(_06145_ ), .A3(_06159_ ), .A4(_06160_ ), .ZN(_00559_ ) );
NOR4_X1 _13747_ ( .A1(_06121_ ), .A2(_04450_ ), .A3(_06144_ ), .A4(_06155_ ), .ZN(_00560_ ) );
NOR4_X1 _13748_ ( .A1(_06121_ ), .A2(\u_lsu.rcount[0] ), .A3(_00879_ ), .A4(_06159_ ), .ZN(_00561_ ) );
AND2_X1 _13749_ ( .A1(\u_lsu.u_clint.mtime[31] ), .A2(\u_lsu.u_clint.mtime[30] ), .ZN(_06161_ ) );
AND2_X1 _13750_ ( .A1(\u_lsu.u_clint.mtime[19] ), .A2(\u_lsu.u_clint.mtime[18] ), .ZN(_06162_ ) );
AND2_X1 _13751_ ( .A1(\u_lsu.u_clint.mtime[17] ), .A2(\u_lsu.u_clint.mtime[16] ), .ZN(_06163_ ) );
AND2_X1 _13752_ ( .A1(_06162_ ), .A2(_06163_ ), .ZN(_06164_ ) );
AND2_X1 _13753_ ( .A1(\u_lsu.u_clint.mtime[23] ), .A2(\u_lsu.u_clint.mtime[22] ), .ZN(_06165_ ) );
AND2_X1 _13754_ ( .A1(\u_lsu.u_clint.mtime[21] ), .A2(\u_lsu.u_clint.mtime[20] ), .ZN(_06166_ ) );
AND3_X1 _13755_ ( .A1(_06164_ ), .A2(_06165_ ), .A3(_06166_ ), .ZN(_06167_ ) );
AND2_X1 _13756_ ( .A1(\u_lsu.u_clint.mtime[29] ), .A2(\u_lsu.u_clint.mtime[28] ), .ZN(_06168_ ) );
AND2_X1 _13757_ ( .A1(\u_lsu.u_clint.mtime[27] ), .A2(\u_lsu.u_clint.mtime[26] ), .ZN(_06169_ ) );
AND2_X1 _13758_ ( .A1(\u_lsu.u_clint.mtime[25] ), .A2(\u_lsu.u_clint.mtime[24] ), .ZN(_06170_ ) );
AND2_X1 _13759_ ( .A1(_06169_ ), .A2(_06170_ ), .ZN(_06171_ ) );
AND4_X1 _13760_ ( .A1(_06161_ ), .A2(_06167_ ), .A3(_06168_ ), .A4(_06171_ ), .ZN(_06172_ ) );
NAND3_X4 _13761_ ( .A1(\u_lsu.u_clint.mtime[1] ), .A2(\u_lsu.u_clint.mtime[2] ), .A3(\u_lsu.u_clint.mtime[0] ), .ZN(_06173_ ) );
NOR2_X2 _13762_ ( .A1(_06173_ ), .A2(_02593_ ), .ZN(_06174_ ) );
AND4_X1 _13763_ ( .A1(\u_lsu.u_clint.mtime[7] ), .A2(\u_lsu.u_clint.mtime[5] ), .A3(\u_lsu.u_clint.mtime[6] ), .A4(\u_lsu.u_clint.mtime[4] ), .ZN(_06175_ ) );
AND2_X1 _13764_ ( .A1(_06174_ ), .A2(_06175_ ), .ZN(_06176_ ) );
INV_X1 _13765_ ( .A(_06176_ ), .ZN(_06177_ ) );
AND2_X1 _13766_ ( .A1(\u_lsu.u_clint.mtime[9] ), .A2(\u_lsu.u_clint.mtime[8] ), .ZN(_06178_ ) );
AND3_X1 _13767_ ( .A1(_06178_ ), .A2(\u_lsu.u_clint.mtime[11] ), .A3(\u_lsu.u_clint.mtime[10] ), .ZN(_06179_ ) );
AND2_X1 _13768_ ( .A1(\u_lsu.u_clint.mtime[15] ), .A2(\u_lsu.u_clint.mtime[14] ), .ZN(_06180_ ) );
NAND4_X1 _13769_ ( .A1(_06179_ ), .A2(\u_lsu.u_clint.mtime[13] ), .A3(\u_lsu.u_clint.mtime[12] ), .A4(_06180_ ), .ZN(_06181_ ) );
NOR2_X1 _13770_ ( .A1(_06177_ ), .A2(_06181_ ), .ZN(_06182_ ) );
AND2_X2 _13771_ ( .A1(_06172_ ), .A2(_06182_ ), .ZN(_06183_ ) );
AND2_X1 _13772_ ( .A1(\u_lsu.u_clint.mtime[35] ), .A2(\u_lsu.u_clint.mtime[34] ), .ZN(_06184_ ) );
AND2_X1 _13773_ ( .A1(\u_lsu.u_clint.mtime[33] ), .A2(\u_lsu.u_clint.mtime[32] ), .ZN(_06185_ ) );
AND2_X1 _13774_ ( .A1(_06184_ ), .A2(_06185_ ), .ZN(_06186_ ) );
AND2_X1 _13775_ ( .A1(\u_lsu.u_clint.mtime[39] ), .A2(\u_lsu.u_clint.mtime[38] ), .ZN(_06187_ ) );
AND2_X1 _13776_ ( .A1(\u_lsu.u_clint.mtime[37] ), .A2(\u_lsu.u_clint.mtime[36] ), .ZN(_06188_ ) );
AND3_X1 _13777_ ( .A1(_06186_ ), .A2(_06187_ ), .A3(_06188_ ), .ZN(_06189_ ) );
AND2_X1 _13778_ ( .A1(\u_lsu.u_clint.mtime[45] ), .A2(\u_lsu.u_clint.mtime[44] ), .ZN(_06190_ ) );
AND3_X1 _13779_ ( .A1(_06190_ ), .A2(\u_lsu.u_clint.mtime[47] ), .A3(\u_lsu.u_clint.mtime[46] ), .ZN(_06191_ ) );
AND2_X1 _13780_ ( .A1(\u_lsu.u_clint.mtime[43] ), .A2(\u_lsu.u_clint.mtime[42] ), .ZN(_06192_ ) );
AND2_X1 _13781_ ( .A1(\u_lsu.u_clint.mtime[41] ), .A2(\u_lsu.u_clint.mtime[40] ), .ZN(_06193_ ) );
AND2_X1 _13782_ ( .A1(_06192_ ), .A2(_06193_ ), .ZN(_06194_ ) );
AND3_X1 _13783_ ( .A1(_06189_ ), .A2(_06191_ ), .A3(_06194_ ), .ZN(_06195_ ) );
AND2_X1 _13784_ ( .A1(_06183_ ), .A2(_06195_ ), .ZN(_06196_ ) );
AND2_X1 _13785_ ( .A1(\u_lsu.u_clint.mtime[51] ), .A2(\u_lsu.u_clint.mtime[50] ), .ZN(_06197_ ) );
AND2_X1 _13786_ ( .A1(\u_lsu.u_clint.mtime[49] ), .A2(\u_lsu.u_clint.mtime[48] ), .ZN(_06198_ ) );
AND2_X1 _13787_ ( .A1(_06197_ ), .A2(_06198_ ), .ZN(_06199_ ) );
AND2_X1 _13788_ ( .A1(\u_lsu.u_clint.mtime[53] ), .A2(\u_lsu.u_clint.mtime[52] ), .ZN(_06200_ ) );
AND4_X1 _13789_ ( .A1(\u_lsu.u_clint.mtime[55] ), .A2(_06199_ ), .A3(\u_lsu.u_clint.mtime[54] ), .A4(_06200_ ), .ZN(_06201_ ) );
AND2_X1 _13790_ ( .A1(_06196_ ), .A2(_06201_ ), .ZN(_06202_ ) );
AND4_X1 _13791_ ( .A1(\u_lsu.u_clint.mtime[59] ), .A2(\u_lsu.u_clint.mtime[57] ), .A3(\u_lsu.u_clint.mtime[58] ), .A4(\u_lsu.u_clint.mtime[56] ), .ZN(_06203_ ) );
AND2_X1 _13792_ ( .A1(_06202_ ), .A2(_06203_ ), .ZN(_06204_ ) );
AND3_X1 _13793_ ( .A1(_06204_ ), .A2(\u_lsu.u_clint.mtime[61] ), .A3(\u_lsu.u_clint.mtime[60] ), .ZN(_06205_ ) );
INV_X1 _13794_ ( .A(_06205_ ), .ZN(_06206_ ) );
OR3_X1 _13795_ ( .A1(_06206_ ), .A2(\u_lsu.u_clint.mtime[63] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ), .ZN(_06207_ ) );
OAI21_X1 _13796_ ( .A(\u_lsu.u_clint.mtime[63] ), .B1(_06206_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ), .ZN(_06208_ ) );
AOI21_X1 _13797_ ( .A(_04454_ ), .B1(_06207_ ), .B2(_06208_ ), .ZN(_00562_ ) );
XNOR2_X1 _13798_ ( .A(_06205_ ), .B(\u_lsu.u_clint.mtime[62] ), .ZN(_06209_ ) );
NOR2_X1 _13799_ ( .A1(_06209_ ), .A2(_04475_ ), .ZN(_00563_ ) );
AND2_X1 _13800_ ( .A1(\u_lsu.u_clint.mtime[5] ), .A2(\u_lsu.u_clint.mtime[4] ), .ZN(_06210_ ) );
AND2_X4 _13801_ ( .A1(_06174_ ), .A2(_06210_ ), .ZN(_06211_ ) );
NAND4_X1 _13802_ ( .A1(_06211_ ), .A2(\u_lsu.u_clint.mtime[7] ), .A3(\u_lsu.u_clint.mtime[9] ), .A4(\u_lsu.u_clint.mtime[6] ), .ZN(_06212_ ) );
INV_X1 _13803_ ( .A(\u_lsu.u_clint.mtime[8] ), .ZN(_06213_ ) );
NOR2_X1 _13804_ ( .A1(_06212_ ), .A2(_06213_ ), .ZN(_06214_ ) );
AND4_X1 _13805_ ( .A1(\u_lsu.u_clint.mtime[13] ), .A2(_06214_ ), .A3(\u_lsu.u_clint.mtime[11] ), .A4(\u_lsu.u_clint.mtime[10] ), .ZN(_06215_ ) );
AND3_X1 _13806_ ( .A1(_06215_ ), .A2(\u_lsu.u_clint.mtime[15] ), .A3(\u_lsu.u_clint.mtime[12] ), .ZN(_06216_ ) );
NAND2_X1 _13807_ ( .A1(_06216_ ), .A2(\u_lsu.u_clint.mtime[14] ), .ZN(_06217_ ) );
INV_X1 _13808_ ( .A(\u_lsu.u_clint.mtime[16] ), .ZN(_06218_ ) );
NOR4_X1 _13809_ ( .A1(_06217_ ), .A2(_01725_ ), .A3(_01890_ ), .A4(_06218_ ), .ZN(_06219_ ) );
NAND3_X1 _13810_ ( .A1(_06219_ ), .A2(\u_lsu.u_clint.mtime[21] ), .A3(\u_lsu.u_clint.mtime[18] ), .ZN(_06220_ ) );
INV_X1 _13811_ ( .A(\u_lsu.u_clint.mtime[20] ), .ZN(_06221_ ) );
NOR3_X1 _13812_ ( .A1(_06220_ ), .A2(_01264_ ), .A3(_06221_ ), .ZN(_06222_ ) );
NAND2_X1 _13813_ ( .A1(_06222_ ), .A2(\u_lsu.u_clint.mtime[22] ), .ZN(_06223_ ) );
INV_X1 _13814_ ( .A(\u_lsu.u_clint.mtime[24] ), .ZN(_06224_ ) );
NOR4_X1 _13815_ ( .A1(_06223_ ), .A2(_01730_ ), .A3(_01885_ ), .A4(_06224_ ), .ZN(_06225_ ) );
AND2_X1 _13816_ ( .A1(_06225_ ), .A2(\u_lsu.u_clint.mtime[26] ), .ZN(_06226_ ) );
AND2_X1 _13817_ ( .A1(_06226_ ), .A2(_06168_ ), .ZN(_06227_ ) );
AND2_X1 _13818_ ( .A1(_06227_ ), .A2(_06161_ ), .ZN(_06228_ ) );
AND2_X1 _13819_ ( .A1(_06228_ ), .A2(_06185_ ), .ZN(_06229_ ) );
AND2_X1 _13820_ ( .A1(_06229_ ), .A2(_06184_ ), .ZN(_06230_ ) );
AND2_X1 _13821_ ( .A1(_06230_ ), .A2(_06188_ ), .ZN(_06231_ ) );
AND2_X1 _13822_ ( .A1(_06231_ ), .A2(_06187_ ), .ZN(_06232_ ) );
AND2_X1 _13823_ ( .A1(_06232_ ), .A2(_06193_ ), .ZN(_06233_ ) );
AND2_X1 _13824_ ( .A1(_06233_ ), .A2(_06192_ ), .ZN(_06234_ ) );
NAND2_X1 _13825_ ( .A1(_06234_ ), .A2(_06191_ ), .ZN(_06235_ ) );
INV_X1 _13826_ ( .A(_06198_ ), .ZN(_06236_ ) );
NOR2_X1 _13827_ ( .A1(_06235_ ), .A2(_06236_ ), .ZN(_06237_ ) );
INV_X1 _13828_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_10_A_$_ANDNOT__Y_B ), .ZN(_06238_ ) );
NAND3_X1 _13829_ ( .A1(_06237_ ), .A2(_06238_ ), .A3(_06197_ ), .ZN(_06239_ ) );
INV_X1 _13830_ ( .A(\u_lsu.u_clint.mtime[53] ), .ZN(_06240_ ) );
AOI21_X1 _13831_ ( .A(_01075_ ), .B1(_06239_ ), .B2(_06240_ ), .ZN(_06241_ ) );
AND2_X1 _13832_ ( .A1(\u_lsu.u_clint.mtime[7] ), .A2(\u_lsu.u_clint.mtime[6] ), .ZN(_06242_ ) );
AND3_X1 _13833_ ( .A1(_06211_ ), .A2(_06178_ ), .A3(_06242_ ), .ZN(_06243_ ) );
AND3_X2 _13834_ ( .A1(_06243_ ), .A2(\u_lsu.u_clint.mtime[11] ), .A3(\u_lsu.u_clint.mtime[10] ), .ZN(_06244_ ) );
NAND2_X1 _13835_ ( .A1(_06244_ ), .A2(\u_lsu.u_clint.mtime[12] ), .ZN(_06245_ ) );
INV_X1 _13836_ ( .A(\u_lsu.u_clint.mtime[13] ), .ZN(_06246_ ) );
NOR2_X2 _13837_ ( .A1(_06245_ ), .A2(_06246_ ), .ZN(_06247_ ) );
AND2_X1 _13838_ ( .A1(_06247_ ), .A2(_06180_ ), .ZN(_06248_ ) );
AND2_X4 _13839_ ( .A1(_06248_ ), .A2(_06163_ ), .ZN(_06249_ ) );
AND2_X4 _13840_ ( .A1(_06249_ ), .A2(_06162_ ), .ZN(_06250_ ) );
AND2_X2 _13841_ ( .A1(_06250_ ), .A2(_06166_ ), .ZN(_06251_ ) );
AND2_X4 _13842_ ( .A1(_06251_ ), .A2(_06165_ ), .ZN(_06252_ ) );
AND2_X4 _13843_ ( .A1(_06252_ ), .A2(_06170_ ), .ZN(_06253_ ) );
AND2_X4 _13844_ ( .A1(_06253_ ), .A2(_06169_ ), .ZN(_06254_ ) );
AND2_X1 _13845_ ( .A1(_06254_ ), .A2(_06168_ ), .ZN(_06255_ ) );
AND2_X2 _13846_ ( .A1(_06255_ ), .A2(_06161_ ), .ZN(_06256_ ) );
AND2_X1 _13847_ ( .A1(_06256_ ), .A2(_06185_ ), .ZN(_06257_ ) );
AND2_X1 _13848_ ( .A1(_06257_ ), .A2(_06184_ ), .ZN(_06258_ ) );
AND2_X1 _13849_ ( .A1(_06258_ ), .A2(_06188_ ), .ZN(_06259_ ) );
AND2_X2 _13850_ ( .A1(_06259_ ), .A2(_06187_ ), .ZN(_06260_ ) );
AND2_X4 _13851_ ( .A1(_06260_ ), .A2(_06193_ ), .ZN(_06261_ ) );
AND2_X4 _13852_ ( .A1(_06261_ ), .A2(_06192_ ), .ZN(_06262_ ) );
AND2_X1 _13853_ ( .A1(_06262_ ), .A2(_06191_ ), .ZN(_06263_ ) );
AND2_X2 _13854_ ( .A1(_06263_ ), .A2(_06198_ ), .ZN(_06264_ ) );
NAND4_X1 _13855_ ( .A1(_06264_ ), .A2(\u_lsu.u_clint.mtime[53] ), .A3(_06238_ ), .A4(_06197_ ), .ZN(_06265_ ) );
AND2_X1 _13856_ ( .A1(_06241_ ), .A2(_06265_ ), .ZN(_00564_ ) );
AND2_X1 _13857_ ( .A1(_06196_ ), .A2(_06199_ ), .ZN(_06266_ ) );
XNOR2_X1 _13858_ ( .A(_06266_ ), .B(\u_lsu.u_clint.mtime[52] ), .ZN(_06267_ ) );
NOR2_X1 _13859_ ( .A1(_06267_ ), .A2(_04475_ ), .ZN(_00565_ ) );
NOR3_X1 _13860_ ( .A1(_06235_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ), .A3(_06236_ ), .ZN(_06268_ ) );
OAI21_X1 _13861_ ( .A(_01060_ ), .B1(_06268_ ), .B2(\u_lsu.u_clint.mtime[51] ), .ZN(_06269_ ) );
INV_X1 _13862_ ( .A(_06263_ ), .ZN(_06270_ ) );
NOR3_X1 _13863_ ( .A1(_06270_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ), .A3(_06236_ ), .ZN(_06271_ ) );
AOI21_X1 _13864_ ( .A(_06269_ ), .B1(_06271_ ), .B2(\u_lsu.u_clint.mtime[51] ), .ZN(_00566_ ) );
AND3_X1 _13865_ ( .A1(_06183_ ), .A2(_06198_ ), .A3(_06195_ ), .ZN(_06272_ ) );
XNOR2_X1 _13866_ ( .A(_06272_ ), .B(\u_lsu.u_clint.mtime[50] ), .ZN(_06273_ ) );
NOR2_X1 _13867_ ( .A1(_06273_ ), .A2(_04475_ ), .ZN(_00567_ ) );
NOR2_X1 _13868_ ( .A1(_06235_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ), .ZN(_06274_ ) );
OAI21_X1 _13869_ ( .A(_01060_ ), .B1(_06274_ ), .B2(\u_lsu.u_clint.mtime[49] ), .ZN(_06275_ ) );
INV_X1 _13870_ ( .A(_06262_ ), .ZN(_06276_ ) );
INV_X1 _13871_ ( .A(_06191_ ), .ZN(_06277_ ) );
NOR3_X1 _13872_ ( .A1(_06276_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ), .A3(_06277_ ), .ZN(_06278_ ) );
AOI21_X1 _13873_ ( .A(_06275_ ), .B1(\u_lsu.u_clint.mtime[49] ), .B2(_06278_ ), .ZN(_00568_ ) );
INV_X1 _13874_ ( .A(_06172_ ), .ZN(_06279_ ) );
INV_X1 _13875_ ( .A(_06182_ ), .ZN(_06280_ ) );
INV_X1 _13876_ ( .A(_06195_ ), .ZN(_06281_ ) );
OR4_X1 _13877_ ( .A1(\u_lsu.u_clint.mtime[48] ), .A2(_06279_ ), .A3(_06280_ ), .A4(_06281_ ), .ZN(_06282_ ) );
INV_X1 _13878_ ( .A(_06183_ ), .ZN(_06283_ ) );
OAI21_X1 _13879_ ( .A(\u_lsu.u_clint.mtime[48] ), .B1(_06283_ ), .B2(_06281_ ), .ZN(_06284_ ) );
AOI211_X1 _13880_ ( .A(_00879_ ), .B(_04456_ ), .C1(_06282_ ), .C2(_06284_ ), .ZN(_00569_ ) );
NAND3_X1 _13881_ ( .A1(_06261_ ), .A2(\u_lsu.u_clint.mtime[44] ), .A3(_06192_ ), .ZN(_06285_ ) );
NOR3_X1 _13882_ ( .A1(_06285_ ), .A2(_02115_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ), .ZN(_06286_ ) );
AND2_X1 _13883_ ( .A1(_06286_ ), .A2(\u_lsu.u_clint.mtime[47] ), .ZN(_06287_ ) );
OAI21_X1 _13884_ ( .A(_05410_ ), .B1(_06286_ ), .B2(\u_lsu.u_clint.mtime[47] ), .ZN(_06288_ ) );
NOR2_X1 _13885_ ( .A1(_06287_ ), .A2(_06288_ ), .ZN(_00570_ ) );
AND2_X1 _13886_ ( .A1(_06183_ ), .A2(_06189_ ), .ZN(_06289_ ) );
AND3_X1 _13887_ ( .A1(_06289_ ), .A2(_06190_ ), .A3(_06194_ ), .ZN(_06290_ ) );
XNOR2_X1 _13888_ ( .A(_06290_ ), .B(\u_lsu.u_clint.mtime[46] ), .ZN(_06291_ ) );
NOR2_X1 _13889_ ( .A1(_06291_ ), .A2(_04475_ ), .ZN(_00571_ ) );
INV_X1 _13890_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_18_A_$_ANDNOT__Y_B ), .ZN(_06292_ ) );
NAND3_X1 _13891_ ( .A1(_06261_ ), .A2(_06292_ ), .A3(_06192_ ), .ZN(_06293_ ) );
AOI21_X1 _13892_ ( .A(_01075_ ), .B1(_06293_ ), .B2(_02115_ ), .ZN(_06294_ ) );
NAND4_X1 _13893_ ( .A1(_06261_ ), .A2(\u_lsu.u_clint.mtime[45] ), .A3(_06292_ ), .A4(_06192_ ), .ZN(_06295_ ) );
AND2_X1 _13894_ ( .A1(_06294_ ), .A2(_06295_ ), .ZN(_00572_ ) );
AND2_X1 _13895_ ( .A1(_06289_ ), .A2(_06194_ ), .ZN(_06296_ ) );
XNOR2_X1 _13896_ ( .A(_06296_ ), .B(\u_lsu.u_clint.mtime[44] ), .ZN(_06297_ ) );
NOR2_X1 _13897_ ( .A1(_06297_ ), .A2(_04467_ ), .ZN(_00573_ ) );
INV_X1 _13898_ ( .A(_06204_ ), .ZN(_06298_ ) );
OR3_X1 _13899_ ( .A1(_06298_ ), .A2(\u_lsu.u_clint.mtime[61] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ), .ZN(_06299_ ) );
OAI21_X1 _13900_ ( .A(\u_lsu.u_clint.mtime[61] ), .B1(_06298_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ), .ZN(_06300_ ) );
AOI21_X1 _13901_ ( .A(_00898_ ), .B1(_06299_ ), .B2(_06300_ ), .ZN(_00574_ ) );
NAND3_X1 _13902_ ( .A1(_06183_ ), .A2(_06193_ ), .A3(_06189_ ), .ZN(_06301_ ) );
OR3_X1 _13903_ ( .A1(_06301_ ), .A2(\u_lsu.u_clint.mtime[43] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ), .ZN(_06302_ ) );
OAI21_X1 _13904_ ( .A(\u_lsu.u_clint.mtime[43] ), .B1(_06301_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ), .ZN(_06303_ ) );
AOI21_X1 _13905_ ( .A(_00898_ ), .B1(_06302_ ), .B2(_06303_ ), .ZN(_00575_ ) );
XNOR2_X1 _13906_ ( .A(_06301_ ), .B(\u_lsu.u_clint.mtime[42] ), .ZN(_06304_ ) );
AND2_X1 _13907_ ( .A1(_06304_ ), .A2(_05397_ ), .ZN(_00576_ ) );
INV_X1 _13908_ ( .A(_06289_ ), .ZN(_06305_ ) );
OR3_X1 _13909_ ( .A1(_06305_ ), .A2(\u_lsu.u_clint.mtime[41] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ), .ZN(_06306_ ) );
OAI21_X1 _13910_ ( .A(\u_lsu.u_clint.mtime[41] ), .B1(_06305_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ), .ZN(_06307_ ) );
AOI21_X1 _13911_ ( .A(_00898_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_00577_ ) );
XNOR2_X1 _13912_ ( .A(_06289_ ), .B(\u_lsu.u_clint.mtime[40] ), .ZN(_06308_ ) );
NOR2_X1 _13913_ ( .A1(_06308_ ), .A2(_04467_ ), .ZN(_00578_ ) );
NAND3_X1 _13914_ ( .A1(_06183_ ), .A2(_06188_ ), .A3(_06186_ ), .ZN(_06309_ ) );
OR3_X1 _13915_ ( .A1(_06309_ ), .A2(\u_lsu.u_clint.mtime[39] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ), .ZN(_06310_ ) );
OAI21_X1 _13916_ ( .A(\u_lsu.u_clint.mtime[39] ), .B1(_06309_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ), .ZN(_06311_ ) );
AOI21_X1 _13917_ ( .A(_00898_ ), .B1(_06310_ ), .B2(_06311_ ), .ZN(_00579_ ) );
XNOR2_X1 _13918_ ( .A(_06309_ ), .B(\u_lsu.u_clint.mtime[38] ), .ZN(_06312_ ) );
AND2_X1 _13919_ ( .A1(_06312_ ), .A2(_05397_ ), .ZN(_00580_ ) );
AND3_X1 _13920_ ( .A1(_06257_ ), .A2(_02554_ ), .A3(_06184_ ), .ZN(_06313_ ) );
OAI21_X1 _13921_ ( .A(_05397_ ), .B1(_06313_ ), .B2(\u_lsu.u_clint.mtime[37] ), .ZN(_06314_ ) );
AND4_X1 _13922_ ( .A1(\u_lsu.u_clint.mtime[37] ), .A2(_06257_ ), .A3(_02554_ ), .A4(_06184_ ), .ZN(_06315_ ) );
NOR2_X1 _13923_ ( .A1(_06314_ ), .A2(_06315_ ), .ZN(_00581_ ) );
AND2_X1 _13924_ ( .A1(_06183_ ), .A2(_06186_ ), .ZN(_06316_ ) );
XNOR2_X1 _13925_ ( .A(_06316_ ), .B(\u_lsu.u_clint.mtime[36] ), .ZN(_06317_ ) );
NOR2_X1 _13926_ ( .A1(_06317_ ), .A2(_04467_ ), .ZN(_00582_ ) );
AND3_X1 _13927_ ( .A1(_06256_ ), .A2(_02666_ ), .A3(_06185_ ), .ZN(_06318_ ) );
OAI21_X1 _13928_ ( .A(_05397_ ), .B1(_06318_ ), .B2(\u_lsu.u_clint.mtime[35] ), .ZN(_06319_ ) );
AND4_X1 _13929_ ( .A1(\u_lsu.u_clint.mtime[35] ), .A2(_06256_ ), .A3(_02666_ ), .A4(_06185_ ), .ZN(_06320_ ) );
NOR2_X1 _13930_ ( .A1(_06319_ ), .A2(_06320_ ), .ZN(_00583_ ) );
AND3_X1 _13931_ ( .A1(_06172_ ), .A2(_06185_ ), .A3(_06182_ ), .ZN(_06321_ ) );
XNOR2_X1 _13932_ ( .A(_06321_ ), .B(\u_lsu.u_clint.mtime[34] ), .ZN(_06322_ ) );
NOR3_X1 _13933_ ( .A1(_06322_ ), .A2(_04450_ ), .A3(_04456_ ), .ZN(_00584_ ) );
XNOR2_X1 _13934_ ( .A(_06204_ ), .B(\u_lsu.u_clint.mtime[60] ), .ZN(_06323_ ) );
NOR2_X1 _13935_ ( .A1(_06323_ ), .A2(_04467_ ), .ZN(_00585_ ) );
AND3_X1 _13936_ ( .A1(_06255_ ), .A2(_02800_ ), .A3(_06161_ ), .ZN(_06324_ ) );
OAI21_X1 _13937_ ( .A(_04468_ ), .B1(_06324_ ), .B2(\u_lsu.u_clint.mtime[33] ), .ZN(_06325_ ) );
AND4_X1 _13938_ ( .A1(\u_lsu.u_clint.mtime[33] ), .A2(_06255_ ), .A3(_02800_ ), .A4(_06161_ ), .ZN(_06326_ ) );
NOR2_X1 _13939_ ( .A1(_06325_ ), .A2(_06326_ ), .ZN(_00586_ ) );
XNOR2_X1 _13940_ ( .A(_06183_ ), .B(\u_lsu.u_clint.mtime[32] ), .ZN(_06327_ ) );
NOR3_X1 _13941_ ( .A1(_05478_ ), .A2(_06327_ ), .A3(_06026_ ), .ZN(_00587_ ) );
NAND3_X1 _13942_ ( .A1(_06254_ ), .A2(_01515_ ), .A3(_06168_ ), .ZN(_06328_ ) );
AOI21_X1 _13943_ ( .A(_01075_ ), .B1(_06328_ ), .B2(_01259_ ), .ZN(_06329_ ) );
NAND4_X1 _13944_ ( .A1(_06254_ ), .A2(\u_lsu.u_clint.mtime[31] ), .A3(_01515_ ), .A4(_06168_ ), .ZN(_06330_ ) );
AND2_X1 _13945_ ( .A1(_06329_ ), .A2(_06330_ ), .ZN(_00588_ ) );
AND2_X1 _13946_ ( .A1(_06182_ ), .A2(_06167_ ), .ZN(_06331_ ) );
NAND3_X1 _13947_ ( .A1(_06331_ ), .A2(_06168_ ), .A3(_06171_ ), .ZN(_06332_ ) );
XNOR2_X1 _13948_ ( .A(_06332_ ), .B(\u_lsu.u_clint.mtime[30] ), .ZN(_06333_ ) );
AND3_X1 _13949_ ( .A1(_06333_ ), .A2(_00866_ ), .A3(_05943_ ), .ZN(_00589_ ) );
NAND3_X1 _13950_ ( .A1(_06253_ ), .A2(_01676_ ), .A3(_06169_ ), .ZN(_06334_ ) );
AOI21_X1 _13951_ ( .A(_00897_ ), .B1(_06334_ ), .B2(_01604_ ), .ZN(_06335_ ) );
NAND4_X1 _13952_ ( .A1(_06253_ ), .A2(\u_lsu.u_clint.mtime[29] ), .A3(_01676_ ), .A4(_06169_ ), .ZN(_06336_ ) );
AND2_X1 _13953_ ( .A1(_06335_ ), .A2(_06336_ ), .ZN(_00590_ ) );
AND2_X1 _13954_ ( .A1(_06331_ ), .A2(_06171_ ), .ZN(_06337_ ) );
XNOR2_X1 _13955_ ( .A(_06337_ ), .B(\u_lsu.u_clint.mtime[28] ), .ZN(_06338_ ) );
NOR3_X1 _13956_ ( .A1(_06338_ ), .A2(_04450_ ), .A3(_04456_ ), .ZN(_00591_ ) );
INV_X1 _13957_ ( .A(_06253_ ), .ZN(_06339_ ) );
NOR3_X1 _13958_ ( .A1(_06339_ ), .A2(_01730_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ), .ZN(_06340_ ) );
NOR2_X1 _13959_ ( .A1(_06220_ ), .A2(_06221_ ), .ZN(_06341_ ) );
AND4_X1 _13960_ ( .A1(\u_lsu.u_clint.mtime[23] ), .A2(_06341_ ), .A3(\u_lsu.u_clint.mtime[25] ), .A4(\u_lsu.u_clint.mtime[22] ), .ZN(_06342_ ) );
NAND2_X1 _13961_ ( .A1(_06342_ ), .A2(\u_lsu.u_clint.mtime[24] ), .ZN(_06343_ ) );
NOR2_X1 _13962_ ( .A1(_06343_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ), .ZN(_06344_ ) );
OAI21_X1 _13963_ ( .A(_01061_ ), .B1(_06344_ ), .B2(\u_lsu.u_clint.mtime[27] ), .ZN(_06345_ ) );
NOR2_X1 _13964_ ( .A1(_06340_ ), .A2(_06345_ ), .ZN(_00592_ ) );
AND3_X1 _13965_ ( .A1(_06182_ ), .A2(_06170_ ), .A3(_06167_ ), .ZN(_06346_ ) );
XNOR2_X1 _13966_ ( .A(_06346_ ), .B(\u_lsu.u_clint.mtime[26] ), .ZN(_06347_ ) );
NOR3_X1 _13967_ ( .A1(flush_$_OR__Y_B ), .A2(_06347_ ), .A3(_04450_ ), .ZN(_00593_ ) );
NAND3_X1 _13968_ ( .A1(_06251_ ), .A2(_01954_ ), .A3(_06165_ ), .ZN(_06348_ ) );
AOI21_X1 _13969_ ( .A(_00897_ ), .B1(_06348_ ), .B2(_01885_ ), .ZN(_06349_ ) );
NAND4_X1 _13970_ ( .A1(_06251_ ), .A2(\u_lsu.u_clint.mtime[25] ), .A3(_01954_ ), .A4(_06165_ ), .ZN(_06350_ ) );
AND2_X1 _13971_ ( .A1(_06349_ ), .A2(_06350_ ), .ZN(_00594_ ) );
NAND4_X1 _13972_ ( .A1(_06341_ ), .A2(\u_lsu.u_clint.mtime[23] ), .A3(\u_lsu.u_clint.mtime[24] ), .A4(\u_lsu.u_clint.mtime[22] ), .ZN(_06351_ ) );
NAND2_X1 _13973_ ( .A1(_06351_ ), .A2(_01061_ ), .ZN(_06352_ ) );
AOI21_X1 _13974_ ( .A(_06352_ ), .B1(_06224_ ), .B2(_06223_ ), .ZN(_00595_ ) );
NAND3_X1 _13975_ ( .A1(_06202_ ), .A2(\u_lsu.u_clint.mtime[57] ), .A3(\u_lsu.u_clint.mtime[56] ), .ZN(_06353_ ) );
OR3_X1 _13976_ ( .A1(_06353_ ), .A2(\u_lsu.u_clint.mtime[59] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ), .ZN(_06354_ ) );
OAI21_X1 _13977_ ( .A(\u_lsu.u_clint.mtime[59] ), .B1(_06353_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ), .ZN(_06355_ ) );
AOI21_X1 _13978_ ( .A(_00898_ ), .B1(_06354_ ), .B2(_06355_ ), .ZN(_00596_ ) );
NAND3_X1 _13979_ ( .A1(_06250_ ), .A2(_02062_ ), .A3(_06166_ ), .ZN(_06356_ ) );
AOI21_X1 _13980_ ( .A(_00897_ ), .B1(_06356_ ), .B2(_01264_ ), .ZN(_06357_ ) );
NAND4_X1 _13981_ ( .A1(_06250_ ), .A2(\u_lsu.u_clint.mtime[23] ), .A3(_02062_ ), .A4(_06166_ ), .ZN(_06358_ ) );
AND2_X1 _13982_ ( .A1(_06357_ ), .A2(_06358_ ), .ZN(_00597_ ) );
NAND3_X1 _13983_ ( .A1(_06182_ ), .A2(_06166_ ), .A3(_06164_ ), .ZN(_06359_ ) );
XNOR2_X1 _13984_ ( .A(_06359_ ), .B(\u_lsu.u_clint.mtime[22] ), .ZN(_06360_ ) );
AND3_X1 _13985_ ( .A1(_05943_ ), .A2(_00866_ ), .A3(_06360_ ), .ZN(_00598_ ) );
NAND3_X1 _13986_ ( .A1(_06249_ ), .A2(_01668_ ), .A3(_06162_ ), .ZN(_06361_ ) );
AOI21_X1 _13987_ ( .A(_00897_ ), .B1(_06361_ ), .B2(_01596_ ), .ZN(_06362_ ) );
NAND4_X1 _13988_ ( .A1(_06249_ ), .A2(\u_lsu.u_clint.mtime[21] ), .A3(_01668_ ), .A4(_06162_ ), .ZN(_06363_ ) );
AND2_X1 _13989_ ( .A1(_06362_ ), .A2(_06363_ ), .ZN(_00599_ ) );
NAND3_X1 _13990_ ( .A1(_06219_ ), .A2(\u_lsu.u_clint.mtime[20] ), .A3(\u_lsu.u_clint.mtime[18] ), .ZN(_06364_ ) );
AND2_X1 _13991_ ( .A1(_06364_ ), .A2(_01060_ ), .ZN(_06365_ ) );
AND2_X1 _13992_ ( .A1(_06219_ ), .A2(\u_lsu.u_clint.mtime[18] ), .ZN(_06366_ ) );
OAI21_X1 _13993_ ( .A(_06365_ ), .B1(\u_lsu.u_clint.mtime[20] ), .B2(_06366_ ), .ZN(_06367_ ) );
INV_X1 _13994_ ( .A(_06367_ ), .ZN(_00600_ ) );
INV_X1 _13995_ ( .A(_06249_ ), .ZN(_06368_ ) );
NOR3_X1 _13996_ ( .A1(_06368_ ), .A2(_01725_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ), .ZN(_06369_ ) );
AND3_X1 _13997_ ( .A1(_06216_ ), .A2(\u_lsu.u_clint.mtime[17] ), .A3(\u_lsu.u_clint.mtime[14] ), .ZN(_06370_ ) );
NAND2_X1 _13998_ ( .A1(_06370_ ), .A2(\u_lsu.u_clint.mtime[16] ), .ZN(_06371_ ) );
NOR2_X1 _13999_ ( .A1(_06371_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ), .ZN(_06372_ ) );
OAI21_X1 _14000_ ( .A(_01061_ ), .B1(_06372_ ), .B2(\u_lsu.u_clint.mtime[19] ), .ZN(_06373_ ) );
NOR2_X1 _14001_ ( .A1(_06369_ ), .A2(_06373_ ), .ZN(_00601_ ) );
AND3_X1 _14002_ ( .A1(_06370_ ), .A2(\u_lsu.u_clint.mtime[18] ), .A3(\u_lsu.u_clint.mtime[16] ), .ZN(_06374_ ) );
NOR2_X1 _14003_ ( .A1(_06374_ ), .A2(_01075_ ), .ZN(_06375_ ) );
AND2_X1 _14004_ ( .A1(_06370_ ), .A2(\u_lsu.u_clint.mtime[16] ), .ZN(_06376_ ) );
OAI21_X1 _14005_ ( .A(_06375_ ), .B1(\u_lsu.u_clint.mtime[18] ), .B2(_06376_ ), .ZN(_06377_ ) );
INV_X1 _14006_ ( .A(_06377_ ), .ZN(_00602_ ) );
NAND3_X1 _14007_ ( .A1(_06247_ ), .A2(_01947_ ), .A3(_06180_ ), .ZN(_06378_ ) );
AOI211_X1 _14008_ ( .A(_00856_ ), .B(_00874_ ), .C1(_06378_ ), .C2(_01890_ ), .ZN(_06379_ ) );
NAND4_X1 _14009_ ( .A1(_06247_ ), .A2(\u_lsu.u_clint.mtime[17] ), .A3(_01947_ ), .A4(_06180_ ), .ZN(_06380_ ) );
NAND2_X1 _14010_ ( .A1(_06379_ ), .A2(_06380_ ), .ZN(_06381_ ) );
INV_X1 _14011_ ( .A(_06381_ ), .ZN(_00603_ ) );
AND2_X1 _14012_ ( .A1(_06215_ ), .A2(\u_lsu.u_clint.mtime[12] ), .ZN(_06382_ ) );
NAND4_X1 _14013_ ( .A1(_06382_ ), .A2(\u_lsu.u_clint.mtime[15] ), .A3(\u_lsu.u_clint.mtime[16] ), .A4(\u_lsu.u_clint.mtime[14] ), .ZN(_06383_ ) );
NAND2_X1 _14014_ ( .A1(_06383_ ), .A2(_01061_ ), .ZN(_06384_ ) );
AOI21_X1 _14015_ ( .A(_06384_ ), .B1(_06218_ ), .B2(_06217_ ), .ZN(_00604_ ) );
NOR3_X1 _14016_ ( .A1(_06245_ ), .A2(_06246_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ), .ZN(_06385_ ) );
OAI211_X1 _14017_ ( .A(_05973_ ), .B(_00864_ ), .C1(_06385_ ), .C2(\u_lsu.u_clint.mtime[15] ), .ZN(_06386_ ) );
NOR4_X1 _14018_ ( .A1(_06245_ ), .A2(_01249_ ), .A3(_06246_ ), .A4(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ), .ZN(_06387_ ) );
NOR2_X1 _14019_ ( .A1(_06386_ ), .A2(_06387_ ), .ZN(_00605_ ) );
NAND3_X1 _14020_ ( .A1(_06215_ ), .A2(\u_lsu.u_clint.mtime[14] ), .A3(\u_lsu.u_clint.mtime[12] ), .ZN(_06388_ ) );
AND3_X1 _14021_ ( .A1(_00864_ ), .A2(_05973_ ), .A3(_06388_ ), .ZN(_06389_ ) );
OAI21_X1 _14022_ ( .A(_06389_ ), .B1(\u_lsu.u_clint.mtime[14] ), .B2(_06382_ ), .ZN(_06390_ ) );
INV_X1 _14023_ ( .A(_06390_ ), .ZN(_00606_ ) );
OR2_X1 _14024_ ( .A1(_06353_ ), .A2(\u_lsu.u_clint.mtime[58] ), .ZN(_06391_ ) );
NAND2_X1 _14025_ ( .A1(_06353_ ), .A2(\u_lsu.u_clint.mtime[58] ), .ZN(_06392_ ) );
AOI21_X1 _14026_ ( .A(_00898_ ), .B1(_06391_ ), .B2(_06392_ ), .ZN(_00607_ ) );
NAND2_X1 _14027_ ( .A1(_06243_ ), .A2(\u_lsu.u_clint.mtime[10] ), .ZN(_06393_ ) );
INV_X1 _14028_ ( .A(\u_lsu.u_clint.mtime[11] ), .ZN(_06394_ ) );
NOR3_X1 _14029_ ( .A1(_06393_ ), .A2(_06394_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ), .ZN(_06395_ ) );
OAI211_X1 _14030_ ( .A(_05973_ ), .B(_00864_ ), .C1(\u_lsu.u_clint.mtime[13] ), .C2(_06395_ ), .ZN(_06396_ ) );
NOR4_X1 _14031_ ( .A1(_06393_ ), .A2(_06246_ ), .A3(_06394_ ), .A4(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ), .ZN(_06397_ ) );
OR2_X1 _14032_ ( .A1(_06396_ ), .A2(_06397_ ), .ZN(_06398_ ) );
INV_X1 _14033_ ( .A(_06398_ ), .ZN(_00608_ ) );
NOR2_X1 _14034_ ( .A1(_06244_ ), .A2(\u_lsu.u_clint.mtime[12] ), .ZN(_06399_ ) );
AND4_X1 _14035_ ( .A1(\u_lsu.u_clint.mtime[11] ), .A2(_06214_ ), .A3(\u_lsu.u_clint.mtime[12] ), .A4(\u_lsu.u_clint.mtime[10] ), .ZN(_06400_ ) );
NOR4_X1 _14036_ ( .A1(_06121_ ), .A2(_04450_ ), .A3(_06399_ ), .A4(_06400_ ), .ZN(_00609_ ) );
NOR3_X1 _14037_ ( .A1(_06212_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ), .A3(_06213_ ), .ZN(_06401_ ) );
NOR2_X1 _14038_ ( .A1(_06401_ ), .A2(\u_lsu.u_clint.mtime[11] ), .ZN(_06402_ ) );
NOR4_X1 _14039_ ( .A1(_06212_ ), .A2(_06394_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ), .A4(_06213_ ), .ZN(_06403_ ) );
NOR4_X1 _14040_ ( .A1(_06121_ ), .A2(_04450_ ), .A3(_06402_ ), .A4(_06403_ ), .ZN(_00610_ ) );
OAI21_X1 _14041_ ( .A(_06393_ ), .B1(_06214_ ), .B2(\u_lsu.u_clint.mtime[10] ), .ZN(_06404_ ) );
NOR4_X1 _14042_ ( .A1(_05972_ ), .A2(reset ), .A3(_05971_ ), .A4(_06404_ ), .ZN(_00611_ ) );
OR3_X1 _14043_ ( .A1(_06177_ ), .A2(\u_lsu.u_clint.mtime[9] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ), .ZN(_06405_ ) );
OAI21_X1 _14044_ ( .A(\u_lsu.u_clint.mtime[9] ), .B1(_06177_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ), .ZN(_06406_ ) );
AOI211_X1 _14045_ ( .A(_00879_ ), .B(_00874_ ), .C1(_06405_ ), .C2(_06406_ ), .ZN(_00612_ ) );
XNOR2_X1 _14046_ ( .A(_06176_ ), .B(\u_lsu.u_clint.mtime[8] ), .ZN(_06407_ ) );
NOR4_X1 _14047_ ( .A1(_05972_ ), .A2(reset ), .A3(_05971_ ), .A4(_06407_ ), .ZN(_00613_ ) );
AND3_X1 _14048_ ( .A1(_06174_ ), .A2(_02466_ ), .A3(_06210_ ), .ZN(_06408_ ) );
XNOR2_X1 _14049_ ( .A(_06408_ ), .B(\u_lsu.u_clint.mtime[7] ), .ZN(_06409_ ) );
NOR4_X1 _14050_ ( .A1(_05972_ ), .A2(reset ), .A3(_00859_ ), .A4(_06409_ ), .ZN(_00614_ ) );
XNOR2_X1 _14051_ ( .A(_06211_ ), .B(\u_lsu.u_clint.mtime[6] ), .ZN(_06410_ ) );
NOR4_X1 _14052_ ( .A1(_04455_ ), .A2(reset ), .A3(_00859_ ), .A4(_06410_ ), .ZN(_00615_ ) );
NOR3_X1 _14053_ ( .A1(_06173_ ), .A2(_02593_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ), .ZN(_06411_ ) );
XNOR2_X1 _14054_ ( .A(_06411_ ), .B(\u_lsu.u_clint.mtime[5] ), .ZN(_06412_ ) );
NOR4_X1 _14055_ ( .A1(_04455_ ), .A2(reset ), .A3(_00859_ ), .A4(_06412_ ), .ZN(_00616_ ) );
XNOR2_X1 _14056_ ( .A(_06174_ ), .B(\u_lsu.u_clint.mtime[4] ), .ZN(_06413_ ) );
NOR4_X1 _14057_ ( .A1(_04455_ ), .A2(reset ), .A3(_00859_ ), .A4(_06413_ ), .ZN(_00617_ ) );
INV_X1 _14058_ ( .A(_06202_ ), .ZN(_06414_ ) );
OR3_X1 _14059_ ( .A1(_06414_ ), .A2(\u_lsu.u_clint.mtime[57] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ), .ZN(_06415_ ) );
OAI21_X1 _14060_ ( .A(\u_lsu.u_clint.mtime[57] ), .B1(_06414_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ), .ZN(_06416_ ) );
AOI21_X1 _14061_ ( .A(_00898_ ), .B1(_06415_ ), .B2(_06416_ ), .ZN(_00618_ ) );
NAND3_X1 _14062_ ( .A1(_02668_ ), .A2(\u_lsu.u_clint.mtime[1] ), .A3(\u_lsu.u_clint.mtime[0] ), .ZN(_06417_ ) );
XNOR2_X1 _14063_ ( .A(_06417_ ), .B(_02593_ ), .ZN(_06418_ ) );
NOR4_X1 _14064_ ( .A1(_04455_ ), .A2(reset ), .A3(_00859_ ), .A4(_06418_ ), .ZN(_00619_ ) );
AND2_X1 _14065_ ( .A1(\u_lsu.u_clint.mtime[1] ), .A2(\u_lsu.u_clint.mtime[0] ), .ZN(_06419_ ) );
OR2_X1 _14066_ ( .A1(_06419_ ), .A2(\u_lsu.u_clint.mtime[2] ), .ZN(_06420_ ) );
AND4_X1 _14067_ ( .A1(_05973_ ), .A2(_00864_ ), .A3(_06173_ ), .A4(_06420_ ), .ZN(_00620_ ) );
NOR2_X1 _14068_ ( .A1(\u_lsu.u_clint.mtime[1] ), .A2(\u_lsu.u_clint.mtime[0] ), .ZN(_06421_ ) );
NOR4_X1 _14069_ ( .A1(_06121_ ), .A2(_00879_ ), .A3(_06419_ ), .A4(_06421_ ), .ZN(_00621_ ) );
AND3_X1 _14070_ ( .A1(_05943_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D[0] ), .A3(_05965_ ), .ZN(_00622_ ) );
XNOR2_X1 _14071_ ( .A(_06202_ ), .B(\u_lsu.u_clint.mtime[56] ), .ZN(_06422_ ) );
NOR2_X1 _14072_ ( .A1(_06422_ ), .A2(_04467_ ), .ZN(_00623_ ) );
NAND3_X1 _14073_ ( .A1(_06264_ ), .A2(_06200_ ), .A3(_06197_ ), .ZN(_06423_ ) );
NOR2_X2 _14074_ ( .A1(_06423_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_8_A_$_ANDNOT__Y_B ), .ZN(_06424_ ) );
AND2_X1 _14075_ ( .A1(_06424_ ), .A2(\u_lsu.u_clint.mtime[55] ), .ZN(_06425_ ) );
OAI21_X1 _14076_ ( .A(_01061_ ), .B1(_06424_ ), .B2(\u_lsu.u_clint.mtime[55] ), .ZN(_06426_ ) );
NOR2_X1 _14077_ ( .A1(_06425_ ), .A2(_06426_ ), .ZN(_00624_ ) );
AND3_X1 _14078_ ( .A1(_06196_ ), .A2(_06200_ ), .A3(_06199_ ), .ZN(_06427_ ) );
XNOR2_X1 _14079_ ( .A(_06427_ ), .B(\u_lsu.u_clint.mtime[54] ), .ZN(_06428_ ) );
NOR2_X1 _14080_ ( .A1(_06428_ ), .A2(_04467_ ), .ZN(_00625_ ) );
INV_X1 _14081_ ( .A(\u_lsu.arvalid ), .ZN(_06429_ ) );
NOR4_X1 _14082_ ( .A1(_04455_ ), .A2(reset ), .A3(_00859_ ), .A4(_06429_ ), .ZN(_00626_ ) );
AND4_X1 _14083_ ( .A1(\ea_errtp[0] ), .A2(_00631_ ), .A3(ea_err ), .A4(exu_valid ), .ZN(_00109_ ) );
BUF_X2 _14084_ ( .A(_01195_ ), .Z(\io_master_arburst[0] ) );
NAND2_X1 _14085_ ( .A1(_01152_ ), .A2(_01154_ ), .ZN(\io_master_araddr[22] ) );
NAND2_X1 _14086_ ( .A1(_01157_ ), .A2(_01159_ ), .ZN(\io_master_araddr[21] ) );
NAND2_X1 _14087_ ( .A1(_01151_ ), .A2(_01153_ ), .ZN(\io_master_araddr[17] ) );
NAND2_X1 _14088_ ( .A1(_01156_ ), .A2(_01158_ ), .ZN(\io_master_araddr[18] ) );
NOR2_X1 _14089_ ( .A1(\io_master_arburst[0] ), .A2(_01258_ ), .ZN(\io_master_araddr[2] ) );
AND2_X1 _14090_ ( .A1(_01273_ ), .A2(\u_arbiter.rmask[1] ), .ZN(\io_master_arsize[0] ) );
AOI21_X1 _14091_ ( .A(_06429_ ), .B1(_01666_ ), .B2(_01667_ ), .ZN(io_master_arvalid ) );
NAND2_X1 _14092_ ( .A1(io_master_awready ), .A2(io_master_awvalid ), .ZN(_06430_ ) );
OAI21_X1 _14093_ ( .A(_06430_ ), .B1(_06143_ ), .B2(\u_lsu.writing ), .ZN(\u_lsu.awvalid_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14094_ ( .A(\al_wmask[1] ), .ZN(_06431_ ) );
NOR2_X1 _14095_ ( .A1(_06431_ ), .A2(\al_wmask[0] ), .ZN(\io_master_awsize[0] ) );
AND2_X1 _14096_ ( .A1(\al_wmask[1] ), .A2(\al_wmask[0] ), .ZN(\io_master_awsize[1] ) );
NOR2_X1 _14097_ ( .A1(_06143_ ), .A2(\u_lsu.writing ), .ZN(_06432_ ) );
OR2_X1 _14098_ ( .A1(_06432_ ), .A2(io_master_bvalid ), .ZN(io_master_bvalid_$_OR__B_Y ) );
INV_X1 _14099_ ( .A(\al_wdata[7] ), .ZN(_06433_ ) );
NOR3_X1 _14100_ ( .A1(_06433_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[7] ) );
INV_X1 _14101_ ( .A(\al_wdata[6] ), .ZN(_06434_ ) );
NOR3_X1 _14102_ ( .A1(_06434_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[6] ) );
INV_X1 _14103_ ( .A(\al_wdata[5] ), .ZN(_06435_ ) );
NOR3_X1 _14104_ ( .A1(_06435_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[5] ) );
INV_X1 _14105_ ( .A(\al_wdata[4] ), .ZN(_06436_ ) );
NOR3_X1 _14106_ ( .A1(_06436_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[4] ) );
INV_X1 _14107_ ( .A(\al_wdata[3] ), .ZN(_06437_ ) );
NOR3_X1 _14108_ ( .A1(_06437_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[3] ) );
INV_X1 _14109_ ( .A(\al_wdata[2] ), .ZN(_06438_ ) );
NOR3_X1 _14110_ ( .A1(_06438_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[2] ) );
INV_X1 _14111_ ( .A(\al_wdata[1] ), .ZN(_06439_ ) );
NOR3_X1 _14112_ ( .A1(_06439_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[1] ) );
INV_X1 _14113_ ( .A(\al_wdata[0] ), .ZN(_06440_ ) );
NOR3_X1 _14114_ ( .A1(_06440_ ), .A2(\io_master_awaddr[0] ), .A3(\io_master_awaddr[1] ), .ZN(\io_master_wdata[0] ) );
INV_X1 _14115_ ( .A(\io_master_awaddr[1] ), .ZN(_06441_ ) );
NOR2_X1 _14116_ ( .A1(_06441_ ), .A2(\io_master_awaddr[0] ), .ZN(_06442_ ) );
NOR2_X1 _14117_ ( .A1(\io_master_awaddr[0] ), .A2(\io_master_awaddr[1] ), .ZN(_06443_ ) );
AOI22_X1 _14118_ ( .A1(_06442_ ), .A2(\al_wdata[15] ), .B1(_06443_ ), .B2(\al_wdata[31] ), .ZN(_06444_ ) );
AND2_X1 _14119_ ( .A1(\io_master_awaddr[0] ), .A2(\io_master_awaddr[1] ), .ZN(_06445_ ) );
INV_X1 _14120_ ( .A(_06445_ ), .ZN(_06446_ ) );
INV_X1 _14121_ ( .A(\al_wdata[23] ), .ZN(_06447_ ) );
INV_X1 _14122_ ( .A(\io_master_awaddr[0] ), .ZN(_06448_ ) );
NOR2_X2 _14123_ ( .A1(_06448_ ), .A2(\io_master_awaddr[1] ), .ZN(_06449_ ) );
INV_X1 _14124_ ( .A(_06449_ ), .ZN(_06450_ ) );
OAI221_X1 _14125_ ( .A(_06444_ ), .B1(_06433_ ), .B2(_06446_ ), .C1(_06447_ ), .C2(_06450_ ), .ZN(\io_master_wdata[31] ) );
AOI22_X1 _14126_ ( .A1(_06449_ ), .A2(\al_wdata[22] ), .B1(_06443_ ), .B2(\al_wdata[30] ), .ZN(_06451_ ) );
INV_X1 _14127_ ( .A(\al_wdata[14] ), .ZN(_06452_ ) );
INV_X1 _14128_ ( .A(_06442_ ), .ZN(_06453_ ) );
BUF_X4 _14129_ ( .A(_06453_ ), .Z(_06454_ ) );
OAI221_X1 _14130_ ( .A(_06451_ ), .B1(_06434_ ), .B2(_06446_ ), .C1(_06452_ ), .C2(_06454_ ), .ZN(\io_master_wdata[30] ) );
BUF_X4 _14131_ ( .A(_06448_ ), .Z(_06455_ ) );
BUF_X4 _14132_ ( .A(_06441_ ), .Z(_06456_ ) );
NAND3_X1 _14133_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[21] ), .ZN(_06457_ ) );
INV_X1 _14134_ ( .A(\al_wdata[13] ), .ZN(_06458_ ) );
OAI221_X1 _14135_ ( .A(_06457_ ), .B1(_06450_ ), .B2(_06458_ ), .C1(_06435_ ), .C2(_06454_ ), .ZN(\io_master_wdata[21] ) );
AOI22_X1 _14136_ ( .A1(_06449_ ), .A2(\al_wdata[12] ), .B1(_06443_ ), .B2(\al_wdata[20] ), .ZN(_06459_ ) );
OAI21_X1 _14137_ ( .A(_06459_ ), .B1(_06436_ ), .B2(_06454_ ), .ZN(\io_master_wdata[20] ) );
NAND3_X1 _14138_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[19] ), .ZN(_06460_ ) );
INV_X1 _14139_ ( .A(\al_wdata[11] ), .ZN(_06461_ ) );
OAI221_X1 _14140_ ( .A(_06460_ ), .B1(_06450_ ), .B2(_06461_ ), .C1(_06437_ ), .C2(_06454_ ), .ZN(\io_master_wdata[19] ) );
NAND3_X1 _14141_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[18] ), .ZN(_06462_ ) );
INV_X1 _14142_ ( .A(\al_wdata[10] ), .ZN(_06463_ ) );
OAI221_X1 _14143_ ( .A(_06462_ ), .B1(_06450_ ), .B2(_06463_ ), .C1(_06438_ ), .C2(_06454_ ), .ZN(\io_master_wdata[18] ) );
NAND3_X1 _14144_ ( .A1(_06455_ ), .A2(_06441_ ), .A3(\al_wdata[17] ), .ZN(_06464_ ) );
INV_X1 _14145_ ( .A(\al_wdata[9] ), .ZN(_06465_ ) );
OAI221_X1 _14146_ ( .A(_06464_ ), .B1(_06450_ ), .B2(_06465_ ), .C1(_06439_ ), .C2(_06454_ ), .ZN(\io_master_wdata[17] ) );
AOI22_X1 _14147_ ( .A1(_06449_ ), .A2(\al_wdata[8] ), .B1(_06443_ ), .B2(\al_wdata[16] ), .ZN(_06466_ ) );
OAI21_X1 _14148_ ( .A(_06466_ ), .B1(_06440_ ), .B2(_06454_ ), .ZN(\io_master_wdata[16] ) );
BUF_X4 _14149_ ( .A(_06450_ ), .Z(_06467_ ) );
INV_X1 _14150_ ( .A(\al_wdata[15] ), .ZN(_06468_ ) );
INV_X1 _14151_ ( .A(_06443_ ), .ZN(_06469_ ) );
OAI22_X1 _14152_ ( .A1(_06467_ ), .A2(_06433_ ), .B1(_06468_ ), .B2(_06469_ ), .ZN(\io_master_wdata[15] ) );
OAI22_X1 _14153_ ( .A1(_06467_ ), .A2(_06434_ ), .B1(_06452_ ), .B2(_06469_ ), .ZN(\io_master_wdata[14] ) );
OAI22_X1 _14154_ ( .A1(_06467_ ), .A2(_06435_ ), .B1(_06458_ ), .B2(_06469_ ), .ZN(\io_master_wdata[13] ) );
NAND3_X1 _14155_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[12] ), .ZN(_06470_ ) );
OAI21_X1 _14156_ ( .A(_06470_ ), .B1(_06467_ ), .B2(_06436_ ), .ZN(\io_master_wdata[12] ) );
AOI22_X1 _14157_ ( .A1(_06442_ ), .A2(\al_wdata[13] ), .B1(_06443_ ), .B2(\al_wdata[29] ), .ZN(_06471_ ) );
NAND3_X1 _14158_ ( .A1(_06456_ ), .A2(\al_wdata[21] ), .A3(\io_master_awaddr[0] ), .ZN(_06472_ ) );
OAI211_X1 _14159_ ( .A(_06471_ ), .B(_06472_ ), .C1(_06435_ ), .C2(_06446_ ), .ZN(\io_master_wdata[29] ) );
OAI22_X1 _14160_ ( .A1(_06467_ ), .A2(_06437_ ), .B1(_06461_ ), .B2(_06469_ ), .ZN(\io_master_wdata[11] ) );
OAI22_X1 _14161_ ( .A1(_06467_ ), .A2(_06438_ ), .B1(_06463_ ), .B2(_06469_ ), .ZN(\io_master_wdata[10] ) );
OAI22_X1 _14162_ ( .A1(_06467_ ), .A2(_06439_ ), .B1(_06465_ ), .B2(_06469_ ), .ZN(\io_master_wdata[9] ) );
NAND3_X1 _14163_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[8] ), .ZN(_06473_ ) );
OAI21_X1 _14164_ ( .A(_06473_ ), .B1(_06467_ ), .B2(_06440_ ), .ZN(\io_master_wdata[8] ) );
AOI22_X1 _14165_ ( .A1(\al_wdata[20] ), .A2(_06449_ ), .B1(_06442_ ), .B2(\al_wdata[12] ), .ZN(_06474_ ) );
NAND3_X1 _14166_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[28] ), .ZN(_06475_ ) );
OAI211_X1 _14167_ ( .A(_06474_ ), .B(_06475_ ), .C1(_06436_ ), .C2(_06446_ ), .ZN(\io_master_wdata[28] ) );
AOI22_X1 _14168_ ( .A1(_06449_ ), .A2(\al_wdata[19] ), .B1(_06445_ ), .B2(\al_wdata[3] ), .ZN(_06476_ ) );
NAND3_X1 _14169_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[27] ), .ZN(_06477_ ) );
OAI211_X1 _14170_ ( .A(_06476_ ), .B(_06477_ ), .C1(_06461_ ), .C2(_06454_ ), .ZN(\io_master_wdata[27] ) );
AOI22_X1 _14171_ ( .A1(_06449_ ), .A2(\al_wdata[18] ), .B1(_06443_ ), .B2(\al_wdata[26] ), .ZN(_06478_ ) );
OAI221_X1 _14172_ ( .A(_06478_ ), .B1(_06438_ ), .B2(_06446_ ), .C1(_06463_ ), .C2(_06453_ ), .ZN(\io_master_wdata[26] ) );
AOI22_X1 _14173_ ( .A1(_06449_ ), .A2(\al_wdata[17] ), .B1(_06445_ ), .B2(\al_wdata[1] ), .ZN(_06479_ ) );
NAND3_X1 _14174_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[25] ), .ZN(_06480_ ) );
OAI211_X1 _14175_ ( .A(_06479_ ), .B(_06480_ ), .C1(_06465_ ), .C2(_06454_ ), .ZN(\io_master_wdata[25] ) );
AOI22_X1 _14176_ ( .A1(\al_wdata[16] ), .A2(_06449_ ), .B1(_06442_ ), .B2(\al_wdata[8] ), .ZN(_06481_ ) );
NAND3_X1 _14177_ ( .A1(_06455_ ), .A2(_06456_ ), .A3(\al_wdata[24] ), .ZN(_06482_ ) );
OAI211_X1 _14178_ ( .A(_06481_ ), .B(_06482_ ), .C1(_06440_ ), .C2(_06446_ ), .ZN(\io_master_wdata[24] ) );
NAND3_X1 _14179_ ( .A1(_06448_ ), .A2(\al_wdata[7] ), .A3(\io_master_awaddr[1] ), .ZN(_06483_ ) );
OAI221_X1 _14180_ ( .A(_06483_ ), .B1(_06469_ ), .B2(_06447_ ), .C1(_06467_ ), .C2(_06468_ ), .ZN(\io_master_wdata[23] ) );
NAND3_X1 _14181_ ( .A1(_06448_ ), .A2(_06441_ ), .A3(\al_wdata[22] ), .ZN(_06484_ ) );
OAI221_X1 _14182_ ( .A(_06484_ ), .B1(_06450_ ), .B2(_06452_ ), .C1(_06434_ ), .C2(_06453_ ), .ZN(\io_master_wdata[22] ) );
NAND2_X1 _14183_ ( .A1(io_master_wready ), .A2(io_master_wlast ), .ZN(_06485_ ) );
OAI21_X1 _14184_ ( .A(_06485_ ), .B1(_06143_ ), .B2(\u_lsu.writing ), .ZN(\u_lsu.wlast_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14185_ ( .A(\al_wmask[0] ), .ZN(_06486_ ) );
AND3_X1 _14186_ ( .A1(_06486_ ), .A2(\al_wmask[1] ), .A3(\io_master_awaddr[1] ), .ZN(_06487_ ) );
NOR2_X1 _14187_ ( .A1(_06487_ ), .A2(\io_master_awsize[1] ), .ZN(_06488_ ) );
OAI21_X1 _14188_ ( .A(_06488_ ), .B1(_06486_ ), .B2(_06446_ ), .ZN(\io_master_wstrb[3] ) );
OAI21_X1 _14189_ ( .A(_06488_ ), .B1(_06486_ ), .B2(_06454_ ), .ZN(\io_master_wstrb[2] ) );
NOR3_X1 _14190_ ( .A1(_06431_ ), .A2(\al_wmask[0] ), .A3(\io_master_awaddr[1] ), .ZN(_06489_ ) );
NOR2_X1 _14191_ ( .A1(_06489_ ), .A2(\io_master_awsize[1] ), .ZN(_06490_ ) );
OAI21_X1 _14192_ ( .A(_06490_ ), .B1(_06486_ ), .B2(_06467_ ), .ZN(\io_master_wstrb[1] ) );
OAI21_X1 _14193_ ( .A(_06490_ ), .B1(_06486_ ), .B2(_06469_ ), .ZN(\io_master_wstrb[0] ) );
NAND2_X1 _14194_ ( .A1(_00632_ ), .A2(_00778_ ), .ZN(_06491_ ) );
OAI22_X1 _14195_ ( .A1(_05951_ ), .A2(_01217_ ), .B1(_00764_ ), .B2(_06491_ ), .ZN(\u_arbiter.rvalid_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14196_ ( .A1(\u_lsu.writing ), .A2(io_master_bvalid ), .ZN(_06492_ ) );
OR2_X1 _14197_ ( .A1(_06143_ ), .A2(_06492_ ), .ZN(_06493_ ) );
NAND4_X1 _14198_ ( .A1(_01218_ ), .A2(_06491_ ), .A3(_01220_ ), .A4(_06493_ ), .ZN(\u_arbiter.working_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14199_ ( .A(_06493_ ), .B1(_06491_ ), .B2(\u_exu.eopt[12] ), .ZN(\u_arbiter.wvalid_$_SDFFE_PP0P__Q_E ) );
NOR4_X1 _14200_ ( .A1(_01394_ ), .A2(_01382_ ), .A3(_01412_ ), .A4(_01405_ ), .ZN(_06494_ ) );
OR4_X1 _14201_ ( .A1(ea_err ), .A2(\u_exu.acsrd[6] ), .A3(\u_exu.acsrd[5] ), .A4(\u_exu.acsrd[4] ), .ZN(_06495_ ) );
NOR2_X1 _14202_ ( .A1(_06495_ ), .A2(\u_exu.acsrd[7] ), .ZN(_06496_ ) );
OAI21_X1 _14203_ ( .A(_00797_ ), .B1(_01379_ ), .B2(_01371_ ), .ZN(_06497_ ) );
OAI21_X1 _14204_ ( .A(_00797_ ), .B1(\u_exu.acsrd[11] ), .B2(\u_exu.acsrd[10] ), .ZN(_06498_ ) );
AND2_X1 _14205_ ( .A1(_06497_ ), .A2(_06498_ ), .ZN(_06499_ ) );
NAND3_X1 _14206_ ( .A1(_06494_ ), .A2(_06496_ ), .A3(_06499_ ), .ZN(_06500_ ) );
NOR3_X1 _14207_ ( .A1(_00763_ ), .A2(_01367_ ), .A3(_06500_ ), .ZN(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AOI21_X1 _14208_ ( .A(ea_err ), .B1(_01404_ ), .B2(\u_exu.acsrd[0] ), .ZN(_06501_ ) );
NOR3_X1 _14209_ ( .A1(_01697_ ), .A2(_01394_ ), .A3(_06501_ ), .ZN(_06502_ ) );
NAND3_X1 _14210_ ( .A1(_06496_ ), .A2(_06502_ ), .A3(_06499_ ), .ZN(_06503_ ) );
NOR3_X1 _14211_ ( .A1(_00763_ ), .A2(_01367_ ), .A3(_06503_ ), .ZN(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y ) );
NOR3_X1 _14212_ ( .A1(_01357_ ), .A2(_01359_ ), .A3(_06501_ ), .ZN(_06504_ ) );
NOR4_X1 _14213_ ( .A1(_01394_ ), .A2(_01362_ ), .A3(_01382_ ), .A4(_01385_ ), .ZN(_06505_ ) );
AND4_X1 _14214_ ( .A1(_01368_ ), .A2(_06499_ ), .A3(_06504_ ), .A4(_06505_ ), .ZN(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
MUX2_X1 _14215_ ( .A(\u_exu.exe_start ), .B(_00631_ ), .S(exu_valid ), .Z(\u_exu.exe_end_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14216_ ( .A(_01054_ ), .B1(_01025_ ), .B2(_00763_ ), .ZN(\u_exu.exe_start_$_SDFFE_PP0P__Q_E ) );
AOI211_X1 _14217_ ( .A(_05392_ ), .B(_05407_ ), .C1(_01218_ ), .C2(_01220_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
AOI211_X1 _14218_ ( .A(_05392_ ), .B(_05424_ ), .C1(_01218_ ), .C2(_01220_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
AOI211_X1 _14219_ ( .A(_01231_ ), .B(_05427_ ), .C1(_01218_ ), .C2(_01220_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_Y_$_ANDNOT__B_Y ) );
BUF_X4 _14220_ ( .A(_01205_ ), .Z(_06506_ ) );
NOR2_X1 _14221_ ( .A1(_01296_ ), .A2(_06506_ ), .ZN(\ac_data[31] ) );
NOR2_X1 _14222_ ( .A1(_01525_ ), .A2(_06506_ ), .ZN(\ac_data[30] ) );
NOR2_X1 _14223_ ( .A1(_01610_ ), .A2(_06506_ ), .ZN(\ac_data[21] ) );
NOR2_X1 _14224_ ( .A1(_01684_ ), .A2(_06506_ ), .ZN(\ac_data[20] ) );
NOR2_X1 _14225_ ( .A1(_01736_ ), .A2(_06506_ ), .ZN(\ac_data[19] ) );
NOR2_X1 _14226_ ( .A1(_01822_ ), .A2(_06506_ ), .ZN(\ac_data[18] ) );
NOR2_X1 _14227_ ( .A1(_01897_ ), .A2(_06506_ ), .ZN(\ac_data[17] ) );
NOR2_X1 _14228_ ( .A1(_01962_ ), .A2(_06506_ ), .ZN(\ac_data[16] ) );
NOR2_X1 _14229_ ( .A1(_02022_ ), .A2(_06506_ ), .ZN(\ac_data[15] ) );
NOR2_X1 _14230_ ( .A1(_02075_ ), .A2(_06506_ ), .ZN(\ac_data[14] ) );
BUF_X4 _14231_ ( .A(_01205_ ), .Z(_06507_ ) );
NOR2_X1 _14232_ ( .A1(_02121_ ), .A2(_06507_ ), .ZN(\ac_data[13] ) );
NOR2_X1 _14233_ ( .A1(_02168_ ), .A2(_06507_ ), .ZN(\ac_data[12] ) );
NOR2_X1 _14234_ ( .A1(_02186_ ), .A2(_06507_ ), .ZN(\ac_data[29] ) );
NOR2_X1 _14235_ ( .A1(_02229_ ), .A2(_06507_ ), .ZN(\ac_data[11] ) );
NOR2_X1 _14236_ ( .A1(_02300_ ), .A2(_06507_ ), .ZN(\ac_data[10] ) );
NOR2_X1 _14237_ ( .A1(_02326_ ), .A2(_06507_ ), .ZN(\ac_data[9] ) );
NOR2_X1 _14238_ ( .A1(_02375_ ), .A2(_06507_ ), .ZN(\ac_data[8] ) );
OAI211_X1 _14239_ ( .A(\io_master_arburst[0] ), .B(_02465_ ), .C1(_01286_ ), .C2(_01290_ ), .ZN(_06508_ ) );
INV_X1 _14240_ ( .A(_06508_ ), .ZN(\ac_data[7] ) );
OAI211_X1 _14241_ ( .A(\io_master_arburst[0] ), .B(_02465_ ), .C1(_02471_ ), .C2(_02474_ ), .ZN(_06509_ ) );
INV_X1 _14242_ ( .A(_06509_ ), .ZN(\ac_data[6] ) );
NAND2_X1 _14243_ ( .A1(_02501_ ), .A2(\io_master_arburst[0] ), .ZN(_06510_ ) );
INV_X1 _14244_ ( .A(_06510_ ), .ZN(\ac_data[5] ) );
NAND2_X1 _14245_ ( .A1(_02560_ ), .A2(\io_master_arburst[0] ), .ZN(_06511_ ) );
INV_X1 _14246_ ( .A(_06511_ ), .ZN(\ac_data[4] ) );
NAND2_X1 _14247_ ( .A1(_02598_ ), .A2(\io_master_arburst[0] ), .ZN(_06512_ ) );
INV_X1 _14248_ ( .A(_06512_ ), .ZN(\ac_data[3] ) );
NAND2_X1 _14249_ ( .A1(_02673_ ), .A2(\io_master_arburst[0] ), .ZN(_06513_ ) );
INV_X1 _14250_ ( .A(_06513_ ), .ZN(\ac_data[2] ) );
NOR2_X1 _14251_ ( .A1(_02698_ ), .A2(_06507_ ), .ZN(\ac_data[28] ) );
NAND2_X1 _14252_ ( .A1(_02743_ ), .A2(\io_master_arburst[0] ), .ZN(_06514_ ) );
INV_X1 _14253_ ( .A(_06514_ ), .ZN(\ac_data[1] ) );
OAI211_X1 _14254_ ( .A(\io_master_arburst[0] ), .B(_02465_ ), .C1(_02798_ ), .C2(_02803_ ), .ZN(_06515_ ) );
INV_X1 _14255_ ( .A(_06515_ ), .ZN(\ac_data[0] ) );
NOR2_X1 _14256_ ( .A1(_02851_ ), .A2(_06507_ ), .ZN(\ac_data[27] ) );
NOR2_X1 _14257_ ( .A1(_02890_ ), .A2(_06507_ ), .ZN(\ac_data[26] ) );
NOR2_X1 _14258_ ( .A1(_02928_ ), .A2(_01205_ ), .ZN(\ac_data[25] ) );
NOR2_X1 _14259_ ( .A1(_02948_ ), .A2(_01205_ ), .ZN(\ac_data[24] ) );
NOR2_X1 _14260_ ( .A1(_03006_ ), .A2(_01205_ ), .ZN(\ac_data[23] ) );
NOR2_X1 _14261_ ( .A1(_03044_ ), .A2(_01205_ ), .ZN(\ac_data[22] ) );
OAI21_X1 _14262_ ( .A(_05955_ ), .B1(_05951_ ), .B2(_01205_ ), .ZN(\u_icache.count_$_SDFFE_PP0P__Q_E ) );
AND3_X1 _14263_ ( .A1(_05948_ ), .A2(_05946_ ), .A3(_05945_ ), .ZN(_06516_ ) );
INV_X1 _14264_ ( .A(_06516_ ), .ZN(_06517_ ) );
OAI21_X1 _14265_ ( .A(_06517_ ), .B1(_05952_ ), .B2(_05979_ ), .ZN(\u_icache.ended_$_SDFFE_PP0P__Q_E ) );
OR2_X1 _14266_ ( .A1(_06516_ ), .A2(\u_icache.ended_$_ANDNOT__B_Y ), .ZN(\u_icache.chvalid_$_SDFFE_PP0P__Q_E ) );
OR2_X1 _14267_ ( .A1(_01078_ ), .A2(\u_exu.exe_end_$_ANDNOT__B_Y ), .ZN(\u_exu.alu_p2_$_SDFFE_PP0P__Q_E ) );
OR2_X1 _14268_ ( .A1(_01078_ ), .A2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(\u_idu.decode_ok_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14269_ ( .A(_05959_ ), .B1(_05979_ ), .B2(_05952_ ), .ZN(\u_ifu.inst_ok_$_SDFFE_PP0P__Q_E ) );
OR2_X1 _14270_ ( .A1(_00762_ ), .A2(_00767_ ), .ZN(_06518_ ) );
OAI21_X1 _14271_ ( .A(_06518_ ), .B1(_05979_ ), .B2(_05952_ ), .ZN(\u_ifu.jpc_ok_$_SDFFE_PP0P__Q_E ) );
NOR4_X1 _14272_ ( .A1(_04455_ ), .A2(reset ), .A3(_06089_ ), .A4(_05955_ ), .ZN(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_Y ) );
NOR4_X1 _14273_ ( .A1(_04455_ ), .A2(reset ), .A3(_05469_ ), .A4(_05955_ ), .ZN(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_B_$_ANDNOT__B_Y ) );
OAI21_X1 _14274_ ( .A(_06006_ ), .B1(_06518_ ), .B2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(\u_ifu.pc_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14275_ ( .A(\u_lsu.arvalid ), .B1(_01681_ ), .B2(io_master_arready ), .ZN(_06519_ ) );
NAND2_X1 _14276_ ( .A1(_06519_ ), .A2(_06142_ ), .ZN(\u_lsu.arvalid_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14277_ ( .A(_01215_ ), .ZN(\u_lsu.rvalid ) );
NOR4_X1 _14278_ ( .A1(_05949_ ), .A2(\fc_addr[4] ), .A3(\u_icache.count[1] ), .A4(\u_icache.count_$_NOT__A_Y ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ) );
NOR4_X1 _14279_ ( .A1(_05949_ ), .A2(_05469_ ), .A3(\u_icache.count[1] ), .A4(\u_icache.count[0] ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_1_Y ) );
NOR4_X1 _14280_ ( .A1(_05949_ ), .A2(_05469_ ), .A3(\u_icache.count[1] ), .A4(\u_icache.count_$_NOT__A_Y ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_2_Y ) );
INV_X1 _14281_ ( .A(\u_icache.count[1] ), .ZN(_06520_ ) );
NOR4_X1 _14282_ ( .A1(_05949_ ), .A2(\fc_addr[4] ), .A3(_06520_ ), .A4(\u_icache.count[0] ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _14283_ ( .A1(_05949_ ), .A2(\fc_addr[4] ), .A3(\u_icache.count[1] ), .A4(\u_icache.count[0] ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_4_Y ) );
NOR4_X1 _14284_ ( .A1(_05949_ ), .A2(_05469_ ), .A3(_06520_ ), .A4(\u_icache.count[0] ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_5_Y ) );
NOR4_X1 _14285_ ( .A1(_05949_ ), .A2(_05469_ ), .A3(_06520_ ), .A4(\u_icache.count_$_NOT__A_Y ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_6_Y ) );
NOR4_X1 _14286_ ( .A1(_05949_ ), .A2(\fc_addr[4] ), .A3(_06520_ ), .A4(\u_icache.count_$_NOT__A_Y ), .ZN(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_7_Y ) );
INV_X1 _14287_ ( .A(_06159_ ), .ZN(_06521_ ) );
OAI21_X1 _14288_ ( .A(_06142_ ), .B1(_01215_ ), .B2(_06521_ ), .ZN(\u_lsu.reading_$_SDFFE_PP0P__Q_E ) );
CLKGATE_X1 _14289_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ), .GCK(_06522_ ) );
CLKGATE_X1 _14290_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_Y_$_ANDNOT__B_Y ), .GCK(_06523_ ) );
CLKGATE_X1 _14291_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_06524_ ) );
CLKGATE_X1 _14292_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06525_ ) );
CLKGATE_X1 _14293_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_06526_ ) );
CLKGATE_X1 _14294_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ), .GCK(_06527_ ) );
CLKGATE_X1 _14295_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_2_Y_$_ANDNOT__B_Y ), .GCK(_06528_ ) );
CLKGATE_X1 _14296_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_06529_ ) );
CLKGATE_X1 _14297_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06530_ ) );
CLKGATE_X1 _14298_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ), .GCK(_06531_ ) );
CLKGATE_X1 _14299_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_06532_ ) );
CLKGATE_X1 _14300_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_06533_ ) );
CLKGATE_X1 _14301_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ), .GCK(_06534_ ) );
CLKGATE_X1 _14302_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ), .GCK(_06535_ ) );
CLKGATE_X1 _14303_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ), .GCK(_06536_ ) );
CLKGATE_X1 _14304_ ( .CK(clock ), .E(io_master_bvalid_$_OR__B_Y ), .GCK(_06537_ ) );
CLKGATE_X1 _14305_ ( .CK(clock ), .E(\u_lsu.wlast_$_SDFFE_PP0P__Q_E ), .GCK(_06538_ ) );
CLKGATE_X1 _14306_ ( .CK(clock ), .E(\u_lsu.reading_$_SDFFE_PP0P__Q_E ), .GCK(_06539_ ) );
CLKGATE_X1 _14307_ ( .CK(clock ), .E(\u_lsu.rvalid ), .GCK(_06540_ ) );
CLKGATE_X1 _14308_ ( .CK(clock ), .E(\u_lsu.awvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06541_ ) );
CLKGATE_X1 _14309_ ( .CK(clock ), .E(\u_lsu.arvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06542_ ) );
CLKGATE_X1 _14310_ ( .CK(clock ), .E(\u_ifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_06543_ ) );
CLKGATE_X1 _14311_ ( .CK(clock ), .E(_00000_ ), .GCK(_06544_ ) );
CLKGATE_X1 _14312_ ( .CK(clock ), .E(\u_ifu.jpc_ok_$_SDFFE_PP0P__Q_E ), .GCK(_06545_ ) );
CLKGATE_X1 _14313_ ( .CK(clock ), .E(\u_ifu.inst_ok_$_SDFFE_PP0P__Q_E ), .GCK(_06546_ ) );
CLKGATE_X1 _14314_ ( .CK(clock ), .E(\u_icache.cready_$_ANDNOT__A_Y ), .GCK(_06547_ ) );
CLKGATE_X1 _14315_ ( .CK(clock ), .E(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .GCK(_06548_ ) );
CLKGATE_X1 _14316_ ( .CK(clock ), .E(\u_idu.decode_ok_$_SDFFE_PP0P__Q_E ), .GCK(_06549_ ) );
CLKGATE_X1 _14317_ ( .CK(clock ), .E(\u_icache.ended_$_SDFFE_PP0P__Q_E ), .GCK(_06550_ ) );
CLKGATE_X1 _14318_ ( .CK(clock ), .E(\u_icache.cvalids_$_SDFFE_PP0P__Q_E ), .GCK(_06551_ ) );
CLKGATE_X1 _14319_ ( .CK(clock ), .E(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_B_$_ANDNOT__B_Y ), .GCK(_06552_ ) );
CLKGATE_X1 _14320_ ( .CK(clock ), .E(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_Y ), .GCK(_06553_ ) );
CLKGATE_X1 _14321_ ( .CK(clock ), .E(\u_icache.count_$_SDFFE_PP0P__Q_E ), .GCK(_06554_ ) );
CLKGATE_X1 _14322_ ( .CK(clock ), .E(\u_icache.chvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06555_ ) );
CLKGATE_X1 _14323_ ( .CK(clock ), .E(\u_icache.cready_$_ANDNOT__B_Y_$_OR__B_Y ), .GCK(_06556_ ) );
CLKGATE_X1 _14324_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_6_Y ), .GCK(_06557_ ) );
CLKGATE_X1 _14325_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_5_Y ), .GCK(_06558_ ) );
CLKGATE_X1 _14326_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_2_Y ), .GCK(_06559_ ) );
CLKGATE_X1 _14327_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_1_Y ), .GCK(_06560_ ) );
CLKGATE_X1 _14328_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_7_Y ), .GCK(_06561_ ) );
CLKGATE_X1 _14329_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_3_Y ), .GCK(_06562_ ) );
CLKGATE_X1 _14330_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ), .GCK(_06563_ ) );
CLKGATE_X1 _14331_ ( .CK(clock ), .E(\u_lsu.reading_$_NAND__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_4_Y ), .GCK(_06564_ ) );
CLKGATE_X1 _14332_ ( .CK(clock ), .E(\u_icache.ended_$_ANDNOT__B_Y ), .GCK(_06565_ ) );
CLKGATE_X1 _14333_ ( .CK(clock ), .E(\u_exu.exe_start_$_SDFFE_PP0P__Q_E ), .GCK(_06566_ ) );
CLKGATE_X1 _14334_ ( .CK(clock ), .E(\u_exu.exe_end_$_SDFFE_PP0P__Q_E ), .GCK(_06567_ ) );
CLKGATE_X1 _14335_ ( .CK(clock ), .E(\u_exu.alu_p2_$_SDFFE_PP0P__Q_E ), .GCK(_06568_ ) );
CLKGATE_X1 _14336_ ( .CK(clock ), .E(\u_exu.exe_end_$_ANDNOT__B_Y ), .GCK(_06569_ ) );
CLKGATE_X1 _14337_ ( .CK(clock ), .E(flush_$_OR__Y_B ), .GCK(_06570_ ) );
CLKGATE_X1 _14338_ ( .CK(clock ), .E(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06571_ ) );
CLKGATE_X1 _14339_ ( .CK(clock ), .E(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y ), .GCK(_06572_ ) );
CLKGATE_X1 _14340_ ( .CK(clock ), .E(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_06573_ ) );
CLKGATE_X1 _14341_ ( .CK(clock ), .E(\u_arbiter.wvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06574_ ) );
CLKGATE_X1 _14342_ ( .CK(clock ), .E(\u_arbiter.working_$_SDFFE_PP0P__Q_E ), .GCK(_06575_ ) );
CLKGATE_X1 _14343_ ( .CK(clock ), .E(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_06576_ ) );
CLKGATE_X1 _14344_ ( .CK(clock ), .E(\u_arbiter.rvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06577_ ) );
CLKGATE_X1 _14345_ ( .CK(clock ), .E(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_AND__A_Y ), .GCK(_06578_ ) );
LOGIC1_X1 _14346_ ( .Z(io_master_bready ) );
LOGIC0_X1 _14347_ ( .Z(\io_master_arburst[1] ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q ( .D(_00001_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[31] ), .QN(_07229_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_1 ( .D(_00002_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[30] ), .QN(_07228_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_10 ( .D(_00003_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[21] ), .QN(_07227_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_11 ( .D(_00004_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[20] ), .QN(_07226_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_12 ( .D(_00005_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[19] ), .QN(_07225_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_13 ( .D(_00006_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[18] ), .QN(_07224_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_14 ( .D(_00007_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[17] ), .QN(_07223_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_15 ( .D(_00008_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[16] ), .QN(_07222_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_16 ( .D(_00009_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[15] ), .QN(_07221_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_17 ( .D(_00010_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[14] ), .QN(_07220_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_18 ( .D(_00011_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[13] ), .QN(_07219_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_19 ( .D(_00012_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[12] ), .QN(_07218_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_2 ( .D(_00013_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[29] ), .QN(_07217_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_20 ( .D(_00014_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[11] ), .QN(_07216_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_21 ( .D(_00015_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[10] ), .QN(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_B ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_22 ( .D(_00016_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[9] ), .QN(_07215_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_23 ( .D(_00017_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[8] ), .QN(io_master_rready_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_24 ( .D(_00018_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[7] ), .QN(_07214_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_25 ( .D(_00019_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[6] ), .QN(io_master_araddr_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_26 ( .D(_00020_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[5] ), .QN(_07213_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_27 ( .D(_00021_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[4] ), .QN(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_B ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_28 ( .D(_00022_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[3] ), .QN(_07212_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_29 ( .D(_00023_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[2] ), .QN(_07211_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_3 ( .D(_00024_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[28] ), .QN(_07210_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_30 ( .D(_00025_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[1] ), .QN(_07209_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_31 ( .D(_00026_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[0] ), .QN(_07208_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_4 ( .D(_00027_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[27] ), .QN(_07207_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_5 ( .D(_00028_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[26] ), .QN(_07206_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_6 ( .D(_00029_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[25] ), .QN(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_B ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_7 ( .D(_00030_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[24] ), .QN(_07205_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_8 ( .D(_00031_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[23] ), .QN(_07204_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_9 ( .D(_00032_ ), .CK(_06578_ ), .Q(\u_arbiter.raddr[22] ), .QN(_07203_ ) );
DFF_X1 \u_arbiter.rmask_$_SDFFE_PP0P__Q ( .D(_00033_ ), .CK(_06578_ ), .Q(\u_arbiter.rmask[1] ), .QN(_07202_ ) );
DFF_X1 \u_arbiter.rmask_$_SDFFE_PP0P__Q_1 ( .D(_00034_ ), .CK(_06578_ ), .Q(\u_arbiter.rmask[0] ), .QN(_07201_ ) );
DFF_X1 \u_arbiter.rsign_$_SDFFE_PP0P__Q ( .D(_00035_ ), .CK(_06578_ ), .Q(\u_arbiter.rsign ), .QN(_07200_ ) );
DFF_X1 \u_arbiter.rvalid_$_SDFFE_PP0P__Q ( .D(_00036_ ), .CK(_06577_ ), .Q(\u_arbiter.rvalid ), .QN(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_A ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q ( .D(_00001_ ), .CK(_06576_ ), .Q(\io_master_awaddr[31] ), .QN(_07199_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_1 ( .D(_00002_ ), .CK(_06576_ ), .Q(\io_master_awaddr[30] ), .QN(_07198_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_10 ( .D(_00003_ ), .CK(_06576_ ), .Q(\io_master_awaddr[21] ), .QN(_07197_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_11 ( .D(_00004_ ), .CK(_06576_ ), .Q(\io_master_awaddr[20] ), .QN(_07196_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_12 ( .D(_00005_ ), .CK(_06576_ ), .Q(\io_master_awaddr[19] ), .QN(_07195_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_13 ( .D(_00006_ ), .CK(_06576_ ), .Q(\io_master_awaddr[18] ), .QN(_07194_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_14 ( .D(_00007_ ), .CK(_06576_ ), .Q(\io_master_awaddr[17] ), .QN(_07193_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_15 ( .D(_00008_ ), .CK(_06576_ ), .Q(\io_master_awaddr[16] ), .QN(_07192_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_16 ( .D(_00009_ ), .CK(_06576_ ), .Q(\io_master_awaddr[15] ), .QN(_07191_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_17 ( .D(_00010_ ), .CK(_06576_ ), .Q(\io_master_awaddr[14] ), .QN(_07190_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_18 ( .D(_00011_ ), .CK(_06576_ ), .Q(\io_master_awaddr[13] ), .QN(_07189_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_19 ( .D(_00012_ ), .CK(_06576_ ), .Q(\io_master_awaddr[12] ), .QN(_07188_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_2 ( .D(_00013_ ), .CK(_06576_ ), .Q(\io_master_awaddr[29] ), .QN(_07187_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_20 ( .D(_00014_ ), .CK(_06576_ ), .Q(\io_master_awaddr[11] ), .QN(_07186_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_21 ( .D(_00015_ ), .CK(_06576_ ), .Q(\io_master_awaddr[10] ), .QN(_07185_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_22 ( .D(_00016_ ), .CK(_06576_ ), .Q(\io_master_awaddr[9] ), .QN(_07184_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_23 ( .D(_00017_ ), .CK(_06576_ ), .Q(\io_master_awaddr[8] ), .QN(_07183_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_24 ( .D(_00018_ ), .CK(_06576_ ), .Q(\io_master_awaddr[7] ), .QN(_07182_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_25 ( .D(_00019_ ), .CK(_06576_ ), .Q(\io_master_awaddr[6] ), .QN(_07181_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_26 ( .D(_00020_ ), .CK(_06576_ ), .Q(\io_master_awaddr[5] ), .QN(_07180_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_27 ( .D(_00021_ ), .CK(_06576_ ), .Q(\io_master_awaddr[4] ), .QN(_07179_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_28 ( .D(_00022_ ), .CK(_06576_ ), .Q(\io_master_awaddr[3] ), .QN(_07178_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_29 ( .D(_00023_ ), .CK(_06576_ ), .Q(\io_master_awaddr[2] ), .QN(_07177_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_3 ( .D(_00024_ ), .CK(_06576_ ), .Q(\io_master_awaddr[28] ), .QN(_07176_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_30 ( .D(_00025_ ), .CK(_06576_ ), .Q(\io_master_awaddr[1] ), .QN(_07175_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_31 ( .D(_00026_ ), .CK(_06576_ ), .Q(\io_master_awaddr[0] ), .QN(_07174_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_4 ( .D(_00027_ ), .CK(_06576_ ), .Q(\io_master_awaddr[27] ), .QN(_07173_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_5 ( .D(_00028_ ), .CK(_06576_ ), .Q(\io_master_awaddr[26] ), .QN(_07172_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_6 ( .D(_00029_ ), .CK(_06576_ ), .Q(\io_master_awaddr[25] ), .QN(_07171_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_7 ( .D(_00030_ ), .CK(_06576_ ), .Q(\io_master_awaddr[24] ), .QN(_07170_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_8 ( .D(_00031_ ), .CK(_06576_ ), .Q(\io_master_awaddr[23] ), .QN(_07169_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_9 ( .D(_00032_ ), .CK(_06576_ ), .Q(\io_master_awaddr[22] ), .QN(_07168_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q ( .D(_00037_ ), .CK(_06578_ ), .Q(\u_arbiter.wbaddr[3] ), .QN(_07167_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q_1 ( .D(_00038_ ), .CK(_06578_ ), .Q(\u_arbiter.wbaddr[2] ), .QN(_07166_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q_2 ( .D(_00039_ ), .CK(_06578_ ), .Q(\u_arbiter.wbaddr[1] ), .QN(_07165_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q_3 ( .D(_00040_ ), .CK(_06578_ ), .Q(\u_arbiter.wbaddr[0] ), .QN(_07164_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q ( .D(_00041_ ), .CK(_06576_ ), .Q(\al_wdata[31] ), .QN(_07163_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_1 ( .D(_00042_ ), .CK(_06576_ ), .Q(\al_wdata[30] ), .QN(_07162_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_10 ( .D(_00043_ ), .CK(_06576_ ), .Q(\al_wdata[21] ), .QN(_07161_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_11 ( .D(_00044_ ), .CK(_06576_ ), .Q(\al_wdata[20] ), .QN(_07160_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_12 ( .D(_00045_ ), .CK(_06576_ ), .Q(\al_wdata[19] ), .QN(_07159_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_13 ( .D(_00046_ ), .CK(_06576_ ), .Q(\al_wdata[18] ), .QN(_07158_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_14 ( .D(_00047_ ), .CK(_06576_ ), .Q(\al_wdata[17] ), .QN(_07157_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_15 ( .D(_00048_ ), .CK(_06576_ ), .Q(\al_wdata[16] ), .QN(_07156_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_16 ( .D(_00049_ ), .CK(_06576_ ), .Q(\al_wdata[15] ), .QN(_07155_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_17 ( .D(_00050_ ), .CK(_06576_ ), .Q(\al_wdata[14] ), .QN(_07154_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_18 ( .D(_00051_ ), .CK(_06576_ ), .Q(\al_wdata[13] ), .QN(_07153_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_19 ( .D(_00052_ ), .CK(_06576_ ), .Q(\al_wdata[12] ), .QN(_07152_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_2 ( .D(_00053_ ), .CK(_06576_ ), .Q(\al_wdata[29] ), .QN(_07151_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_20 ( .D(_00054_ ), .CK(_06576_ ), .Q(\al_wdata[11] ), .QN(_07150_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_21 ( .D(_00055_ ), .CK(_06576_ ), .Q(\al_wdata[10] ), .QN(_07149_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_22 ( .D(_00056_ ), .CK(_06576_ ), .Q(\al_wdata[9] ), .QN(_07148_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_23 ( .D(_00057_ ), .CK(_06576_ ), .Q(\al_wdata[8] ), .QN(_07147_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_24 ( .D(_00058_ ), .CK(_06576_ ), .Q(\al_wdata[7] ), .QN(_07146_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_25 ( .D(_00059_ ), .CK(_06576_ ), .Q(\al_wdata[6] ), .QN(_07145_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_26 ( .D(_00060_ ), .CK(_06576_ ), .Q(\al_wdata[5] ), .QN(_07144_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_27 ( .D(_00061_ ), .CK(_06576_ ), .Q(\al_wdata[4] ), .QN(_07143_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_28 ( .D(_00062_ ), .CK(_06576_ ), .Q(\al_wdata[3] ), .QN(_07142_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_29 ( .D(_00063_ ), .CK(_06576_ ), .Q(\al_wdata[2] ), .QN(_07141_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_3 ( .D(_00064_ ), .CK(_06576_ ), .Q(\al_wdata[28] ), .QN(_07140_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_30 ( .D(_00065_ ), .CK(_06576_ ), .Q(\al_wdata[1] ), .QN(_07139_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_31 ( .D(_00066_ ), .CK(_06576_ ), .Q(\al_wdata[0] ), .QN(_07138_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_4 ( .D(_00067_ ), .CK(_06576_ ), .Q(\al_wdata[27] ), .QN(_07137_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_5 ( .D(_00068_ ), .CK(_06576_ ), .Q(\al_wdata[26] ), .QN(_07136_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_6 ( .D(_00069_ ), .CK(_06576_ ), .Q(\al_wdata[25] ), .QN(_07135_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_7 ( .D(_00070_ ), .CK(_06576_ ), .Q(\al_wdata[24] ), .QN(_07134_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_8 ( .D(_00071_ ), .CK(_06576_ ), .Q(\al_wdata[23] ), .QN(_07133_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_9 ( .D(_00072_ ), .CK(_06576_ ), .Q(\al_wdata[22] ), .QN(_07132_ ) );
DFF_X1 \u_arbiter.wmask_$_SDFFE_PP0P__Q ( .D(_00033_ ), .CK(_06576_ ), .Q(\al_wmask[1] ), .QN(_07131_ ) );
DFF_X1 \u_arbiter.wmask_$_SDFFE_PP0P__Q_1 ( .D(_00034_ ), .CK(_06576_ ), .Q(\al_wmask[0] ), .QN(_07130_ ) );
DFF_X1 \u_arbiter.working_$_SDFFE_PP0P__Q ( .D(_00073_ ), .CK(_06575_ ), .Q(\u_arbiter.working ), .QN(_07129_ ) );
DFF_X1 \u_arbiter.wvalid_$_SDFFE_PP0P__Q ( .D(_00074_ ), .CK(_06574_ ), .Q(\u_arbiter.wvalid ), .QN(_07128_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q ( .D(_00075_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][31] ), .QN(_07127_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_1 ( .D(_00076_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][30] ), .QN(_07126_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_10 ( .D(_00077_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][21] ), .QN(_07125_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_11 ( .D(_00078_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][20] ), .QN(_07124_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_12 ( .D(_00079_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][19] ), .QN(_07123_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_13 ( .D(_00080_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][18] ), .QN(_07122_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_14 ( .D(_00081_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][17] ), .QN(_07121_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_15 ( .D(_00082_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][16] ), .QN(_07120_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_16 ( .D(_00083_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][15] ), .QN(_07119_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_17 ( .D(_00084_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][14] ), .QN(_07118_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_18 ( .D(_00085_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][13] ), .QN(_07117_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_19 ( .D(_00086_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][10] ), .QN(_07116_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_2 ( .D(_00087_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][29] ), .QN(_07115_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_20 ( .D(_00088_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][9] ), .QN(_07114_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_21 ( .D(_00089_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][8] ), .QN(_07113_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_22 ( .D(_00090_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][7] ), .QN(_07112_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_23 ( .D(_00091_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][6] ), .QN(_07111_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_24 ( .D(_00092_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][5] ), .QN(_07110_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_25 ( .D(_00093_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][4] ), .QN(_07109_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_26 ( .D(_00094_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][3] ), .QN(_07108_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_27 ( .D(_00095_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][2] ), .QN(_07107_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_28 ( .D(_00096_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][1] ), .QN(_07106_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_29 ( .D(_00097_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][0] ), .QN(_07105_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_3 ( .D(_00098_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][28] ), .QN(_07104_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_4 ( .D(_00099_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][27] ), .QN(_07103_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_5 ( .D(_00100_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][26] ), .QN(_07102_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_6 ( .D(_00101_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][25] ), .QN(_07101_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_7 ( .D(_00102_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][24] ), .QN(_07100_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_8 ( .D(_00103_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][23] ), .QN(_07099_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_9 ( .D(_00104_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][22] ), .QN(_07098_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP1P__Q ( .D(_00105_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][12] ), .QN(_07097_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP1P__Q_1 ( .D(_00106_ ), .CK(_06573_ ), .Q(\u_csr.csr[0][11] ), .QN(_07096_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q ( .D(_00075_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][31] ), .QN(_07095_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_1 ( .D(_00076_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][30] ), .QN(_07094_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_10 ( .D(_00077_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][21] ), .QN(_07093_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_11 ( .D(_00078_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][20] ), .QN(_07092_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_12 ( .D(_00079_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][19] ), .QN(_07091_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_13 ( .D(_00080_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][18] ), .QN(_07090_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_14 ( .D(_00081_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][17] ), .QN(_07089_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_15 ( .D(_00082_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][16] ), .QN(_07088_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_16 ( .D(_00083_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][15] ), .QN(_07087_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_17 ( .D(_00084_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][14] ), .QN(_07086_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_18 ( .D(_00085_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][13] ), .QN(_07085_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_19 ( .D(_00107_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][12] ), .QN(_07084_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_2 ( .D(_00087_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][29] ), .QN(_07083_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_20 ( .D(_00108_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][11] ), .QN(_07082_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_21 ( .D(_00086_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][10] ), .QN(_07081_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_22 ( .D(_00088_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][9] ), .QN(_07080_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_23 ( .D(_00089_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][8] ), .QN(_07079_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_24 ( .D(_00090_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][7] ), .QN(_07078_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_25 ( .D(_00091_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][6] ), .QN(_07077_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_26 ( .D(_00092_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][5] ), .QN(_07076_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_27 ( .D(_00093_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][4] ), .QN(_07075_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_28 ( .D(_00094_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][3] ), .QN(_07074_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_29 ( .D(_00095_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][2] ), .QN(_07073_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_3 ( .D(_00098_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][28] ), .QN(_07072_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_30 ( .D(_00096_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][1] ), .QN(_07071_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_31 ( .D(_00097_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][0] ), .QN(_07070_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_4 ( .D(_00099_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][27] ), .QN(_07069_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_5 ( .D(_00100_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][26] ), .QN(_07068_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_6 ( .D(_00101_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][25] ), .QN(_07067_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_7 ( .D(_00102_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][24] ), .QN(_07066_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_8 ( .D(_00103_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][23] ), .QN(_07065_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_9 ( .D(_00104_ ), .CK(_06572_ ), .Q(\u_csr.csr[1][22] ), .QN(_07064_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q ( .D(_00075_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][31] ), .QN(_07063_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_1 ( .D(_00076_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][30] ), .QN(_07062_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_10 ( .D(_00077_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][21] ), .QN(_07061_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_11 ( .D(_00078_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][20] ), .QN(_07060_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_12 ( .D(_00079_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][19] ), .QN(_07059_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_13 ( .D(_00080_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][18] ), .QN(_07058_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_14 ( .D(_00081_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][17] ), .QN(_07057_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_15 ( .D(_00082_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][16] ), .QN(_07056_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_16 ( .D(_00083_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][15] ), .QN(_07055_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_17 ( .D(_00084_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][14] ), .QN(_07054_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_18 ( .D(_00085_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][13] ), .QN(_07053_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_19 ( .D(_00107_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][12] ), .QN(_07052_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_2 ( .D(_00087_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][29] ), .QN(_07051_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_20 ( .D(_00108_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][11] ), .QN(_07050_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_21 ( .D(_00086_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][10] ), .QN(_07049_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_22 ( .D(_00088_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][9] ), .QN(_07048_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_23 ( .D(_00089_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][8] ), .QN(_07047_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_24 ( .D(_00090_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][7] ), .QN(_07046_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_25 ( .D(_00091_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][6] ), .QN(_07045_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_26 ( .D(_00092_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][5] ), .QN(_07044_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_27 ( .D(_00093_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][4] ), .QN(_07043_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_28 ( .D(_00094_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][3] ), .QN(_07042_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_29 ( .D(_00095_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][2] ), .QN(_07041_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_3 ( .D(_00098_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][28] ), .QN(_07040_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_30 ( .D(_00096_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][1] ), .QN(_07039_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_31 ( .D(_00097_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][0] ), .QN(_07038_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_4 ( .D(_00099_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][27] ), .QN(_07037_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_5 ( .D(_00100_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][26] ), .QN(_07036_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_6 ( .D(_00101_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][25] ), .QN(_07035_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_7 ( .D(_00102_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][24] ), .QN(_07034_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_8 ( .D(_00103_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][23] ), .QN(_07033_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_9 ( .D(_00104_ ), .CK(_06571_ ), .Q(\u_csr.csr[2][22] ), .QN(_07032_ ) );
DFF_X1 \u_csr.csr[3]_$_SDFFCE_PN0P__Q ( .D(_00109_ ), .CK(_06570_ ), .Q(\u_csr.csr[3][0] ), .QN(_07031_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q ( .D(_00110_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[11] ), .QN(_07030_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_1 ( .D(_00111_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[10] ), .QN(_07029_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_10 ( .D(_00112_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[1] ), .QN(_07028_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_11 ( .D(_00113_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[0] ), .QN(_07027_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_2 ( .D(_00114_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[9] ), .QN(_07026_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_3 ( .D(_00115_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[8] ), .QN(_07025_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_4 ( .D(_00116_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[7] ), .QN(_07024_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_5 ( .D(_00117_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[6] ), .QN(_07023_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_6 ( .D(_00118_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[5] ), .QN(_07022_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_7 ( .D(_00119_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[4] ), .QN(_07021_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_8 ( .D(_00120_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[3] ), .QN(_07020_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_9 ( .D(_00121_ ), .CK(_06569_ ), .Q(\u_exu.acsrd[2] ), .QN(_07019_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q ( .D(_00122_ ), .CK(_06568_ ), .Q(\u_exu.alu_ctrl[6] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_1 ( .D(_00123_ ), .CK(_06568_ ), .Q(\u_exu.alu_ctrl[5] ), .QN(_07018_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_2 ( .D(_00124_ ), .CK(_06568_ ), .Q(\u_exu.alu_ctrl[4] ), .QN(_07017_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_3 ( .D(_00125_ ), .CK(_06568_ ), .Q(\u_exu.alu_ctrl[3] ), .QN(_07016_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_4 ( .D(_00126_ ), .CK(_06568_ ), .Q(\u_exu.alu_ctrl[2] ), .QN(_07015_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_5 ( .D(_00127_ ), .CK(_06568_ ), .Q(\u_exu.alu_ctrl[1] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_Y_$_MUX__B_A_$_NOR__Y_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_6 ( .D(_00128_ ), .CK(_06568_ ), .Q(\u_exu.alu_ctrl[0] ), .QN(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q ( .D(_00129_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[31] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_1 ( .D(_00130_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[30] ), .QN(_07014_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_10 ( .D(_00131_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[21] ), .QN(\u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_11 ( .D(_00132_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[20] ), .QN(_07013_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_12 ( .D(_00133_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[19] ), .QN(\u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_13 ( .D(_00134_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[18] ), .QN(_07012_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_14 ( .D(_00135_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[17] ), .QN(\u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_15 ( .D(_00136_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[16] ), .QN(_07011_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_16 ( .D(_00137_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[15] ), .QN(\u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_17 ( .D(_00138_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[14] ), .QN(_07010_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_18 ( .D(_00139_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[13] ), .QN(_07009_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_19 ( .D(_00140_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[12] ), .QN(_07008_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_2 ( .D(_00141_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[29] ), .QN(_07007_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_20 ( .D(_00142_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[11] ), .QN(\u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_21 ( .D(_00143_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[10] ), .QN(_07006_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_22 ( .D(_00144_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[9] ), .QN(\u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_23 ( .D(_00145_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[8] ), .QN(_07005_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_24 ( .D(_00146_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[7] ), .QN(\u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_25 ( .D(_00147_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[6] ), .QN(_07004_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_26 ( .D(_00148_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[5] ), .QN(\u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_27 ( .D(_00149_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[4] ), .QN(_07003_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_28 ( .D(_00150_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[3] ), .QN(\u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_29 ( .D(_00151_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[2] ), .QN(_07002_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_3 ( .D(_00152_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[28] ), .QN(_07001_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_30 ( .D(_00153_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[1] ), .QN(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_31 ( .D(_00154_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[0] ), .QN(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_4 ( .D(_00155_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[27] ), .QN(_07000_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_5 ( .D(_00156_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[26] ), .QN(_06999_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_6 ( .D(_00157_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[25] ), .QN(_06998_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_7 ( .D(_00158_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[24] ), .QN(_06997_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_8 ( .D(_00159_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[23] ), .QN(_06996_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_9 ( .D(_00160_ ), .CK(_06568_ ), .Q(\u_exu.alu_p1[22] ), .QN(_06995_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q ( .D(_00161_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[31] ), .QN(_06994_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_1 ( .D(_00162_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[30] ), .QN(_06993_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_10 ( .D(_00163_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[21] ), .QN(_06992_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_11 ( .D(_00164_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[20] ), .QN(_06991_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_12 ( .D(_00165_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[19] ), .QN(_06990_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_13 ( .D(_00166_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[18] ), .QN(_06989_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_14 ( .D(_00167_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[17] ), .QN(_06988_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_15 ( .D(_00168_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[16] ), .QN(_06987_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_16 ( .D(_00169_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[15] ), .QN(_06986_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_17 ( .D(_00170_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[14] ), .QN(_06985_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_18 ( .D(_00171_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[13] ), .QN(_06984_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_19 ( .D(_00172_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[12] ), .QN(_06983_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_2 ( .D(_00173_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[29] ), .QN(_06982_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_20 ( .D(_00174_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[11] ), .QN(_06981_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_21 ( .D(_00175_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[10] ), .QN(_06980_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_22 ( .D(_00176_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[9] ), .QN(_06979_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_23 ( .D(_00177_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[8] ), .QN(_06978_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_24 ( .D(_00178_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[7] ), .QN(_06977_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_25 ( .D(_00179_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[6] ), .QN(_06976_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_26 ( .D(_00180_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[5] ), .QN(_06975_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_27 ( .D(_00181_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[4] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B_$_MUX__B_A_$_NAND__Y_B ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_28 ( .D(_00182_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[3] ), .QN(_06974_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_29 ( .D(_00183_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[2] ), .QN(_06973_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_3 ( .D(_00184_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[28] ), .QN(_06972_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_30 ( .D(_00185_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[1] ), .QN(_06971_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_31 ( .D(_00186_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[0] ), .QN(_06970_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_4 ( .D(_00187_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[27] ), .QN(_06969_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_5 ( .D(_00188_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[26] ), .QN(_06968_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_6 ( .D(_00189_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[25] ), .QN(_06967_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_7 ( .D(_00190_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[24] ), .QN(_06966_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_8 ( .D(_00191_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[23] ), .QN(_06965_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_9 ( .D(_00192_ ), .CK(_06568_ ), .Q(\u_exu.alu_p2[22] ), .QN(_06964_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q ( .D(_00193_ ), .CK(_06569_ ), .Q(\ea_ard[3] ), .QN(_06963_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q_1 ( .D(_00194_ ), .CK(_06569_ ), .Q(\ea_ard[2] ), .QN(_06962_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q_2 ( .D(_00195_ ), .CK(_06569_ ), .Q(\ea_ard[1] ), .QN(_06961_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q_3 ( .D(_00196_ ), .CK(_06569_ ), .Q(\ea_ard[0] ), .QN(_06960_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q ( .D(_00197_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[31] ), .QN(_06959_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_1 ( .D(_00198_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[30] ), .QN(_06958_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_10 ( .D(_00199_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[21] ), .QN(_06957_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_11 ( .D(_00200_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[20] ), .QN(_06956_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_12 ( .D(_00201_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[19] ), .QN(_06955_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_13 ( .D(_00202_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[18] ), .QN(_06954_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_14 ( .D(_00203_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[17] ), .QN(_06953_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_15 ( .D(_00204_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[16] ), .QN(_06952_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_16 ( .D(_00205_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[15] ), .QN(_06951_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_17 ( .D(_00206_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[14] ), .QN(_06950_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_18 ( .D(_00207_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[13] ), .QN(_06949_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_19 ( .D(_00208_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[12] ), .QN(_06948_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_2 ( .D(_00209_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[29] ), .QN(_06947_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_20 ( .D(_00210_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[11] ), .QN(_06946_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_21 ( .D(_00211_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[10] ), .QN(_06945_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_22 ( .D(_00212_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[9] ), .QN(_06944_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_23 ( .D(_00213_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[8] ), .QN(_06943_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_24 ( .D(_00214_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[7] ), .QN(_06942_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_25 ( .D(_00215_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[6] ), .QN(_06941_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_26 ( .D(_00216_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[5] ), .QN(_06940_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_27 ( .D(_00217_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[4] ), .QN(_06939_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_28 ( .D(_00218_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[3] ), .QN(_06938_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_29 ( .D(_00219_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[2] ), .QN(_06937_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_3 ( .D(_00220_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[28] ), .QN(_06936_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_30 ( .D(_00221_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[1] ), .QN(_06935_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_31 ( .D(_00222_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[0] ), .QN(_06934_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_4 ( .D(_00223_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[27] ), .QN(_06933_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_5 ( .D(_00224_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[26] ), .QN(_06932_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_6 ( .D(_00225_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[25] ), .QN(_06931_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_7 ( .D(_00226_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[24] ), .QN(_06930_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_8 ( .D(_00227_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[23] ), .QN(_06929_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_9 ( .D(_00228_ ), .CK(_06569_ ), .Q(\u_exu.ecsr[22] ), .QN(_06928_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q ( .D(_00229_ ), .CK(_06569_ ), .Q(\u_exu.eopt[15] ), .QN(_06927_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_1 ( .D(_00230_ ), .CK(_06569_ ), .Q(ea_rsign ), .QN(_06926_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_2 ( .D(_00231_ ), .CK(_06569_ ), .Q(\u_exu.eopt[12] ), .QN(_06925_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_3 ( .D(_00232_ ), .CK(_06569_ ), .Q(\ea_mask[1] ), .QN(_06924_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_4 ( .D(_00233_ ), .CK(_06569_ ), .Q(\ea_mask[0] ), .QN(_06923_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_5 ( .D(_00234_ ), .CK(_06569_ ), .Q(\u_exu.eopt[0] ), .QN(_06922_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q ( .D(_00235_ ), .CK(_06569_ ), .Q(\ea_pc[31] ), .QN(_06921_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_1 ( .D(_00236_ ), .CK(_06569_ ), .Q(\ea_pc[30] ), .QN(_06920_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_10 ( .D(_00237_ ), .CK(_06569_ ), .Q(\ea_pc[21] ), .QN(_06919_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_11 ( .D(_00238_ ), .CK(_06569_ ), .Q(\ea_pc[20] ), .QN(_06918_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_12 ( .D(_00239_ ), .CK(_06569_ ), .Q(\ea_pc[19] ), .QN(_06917_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_13 ( .D(_00240_ ), .CK(_06569_ ), .Q(\ea_pc[18] ), .QN(_06916_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_14 ( .D(_00241_ ), .CK(_06569_ ), .Q(\ea_pc[17] ), .QN(_06915_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_15 ( .D(_00242_ ), .CK(_06569_ ), .Q(\ea_pc[16] ), .QN(_06914_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_16 ( .D(_00243_ ), .CK(_06569_ ), .Q(\ea_pc[15] ), .QN(_06913_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_17 ( .D(_00244_ ), .CK(_06569_ ), .Q(\ea_pc[14] ), .QN(_06912_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_18 ( .D(_00245_ ), .CK(_06569_ ), .Q(\ea_pc[13] ), .QN(_06911_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_19 ( .D(_00246_ ), .CK(_06569_ ), .Q(\ea_pc[12] ), .QN(_06910_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_2 ( .D(_00247_ ), .CK(_06569_ ), .Q(\ea_pc[29] ), .QN(_06909_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_20 ( .D(_00248_ ), .CK(_06569_ ), .Q(\ea_pc[11] ), .QN(_06908_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_21 ( .D(_00249_ ), .CK(_06569_ ), .Q(\ea_pc[10] ), .QN(_06907_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_22 ( .D(_00250_ ), .CK(_06569_ ), .Q(\ea_pc[9] ), .QN(_06906_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_23 ( .D(_00251_ ), .CK(_06569_ ), .Q(\ea_pc[8] ), .QN(_06905_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_24 ( .D(_00252_ ), .CK(_06569_ ), .Q(\ea_pc[7] ), .QN(_06904_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_25 ( .D(_00253_ ), .CK(_06569_ ), .Q(\ea_pc[6] ), .QN(_06903_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_26 ( .D(_00254_ ), .CK(_06569_ ), .Q(\ea_pc[5] ), .QN(_06902_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_27 ( .D(_00255_ ), .CK(_06569_ ), .Q(\ea_pc[4] ), .QN(_06901_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_28 ( .D(_00256_ ), .CK(_06569_ ), .Q(\ea_pc[3] ), .QN(_06900_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_29 ( .D(_00257_ ), .CK(_06569_ ), .Q(\ea_pc[2] ), .QN(_06899_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_3 ( .D(_00258_ ), .CK(_06569_ ), .Q(\ea_pc[28] ), .QN(_06898_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_30 ( .D(_00259_ ), .CK(_06569_ ), .Q(\ea_pc[1] ), .QN(_06897_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_31 ( .D(_00260_ ), .CK(_06569_ ), .Q(\ea_pc[0] ), .QN(_06896_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_4 ( .D(_00261_ ), .CK(_06569_ ), .Q(\ea_pc[27] ), .QN(_06895_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_5 ( .D(_00262_ ), .CK(_06569_ ), .Q(\ea_pc[26] ), .QN(_06894_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_6 ( .D(_00263_ ), .CK(_06569_ ), .Q(\ea_pc[25] ), .QN(_06893_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_7 ( .D(_00264_ ), .CK(_06569_ ), .Q(\ea_pc[24] ), .QN(_06892_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_8 ( .D(_00265_ ), .CK(_06569_ ), .Q(\ea_pc[23] ), .QN(_06891_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_9 ( .D(_00266_ ), .CK(_06569_ ), .Q(\ea_pc[22] ), .QN(_06890_ ) );
DFF_X1 \u_exu.error_$_SDFFE_PP0P__Q ( .D(_00267_ ), .CK(_06569_ ), .Q(ea_err ), .QN(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ) );
DFF_X1 \u_exu.errtp_$_SDFFE_PP0P__Q ( .D(_00268_ ), .CK(_06569_ ), .Q(\ea_errtp[0] ), .QN(_06889_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q ( .D(_00269_ ), .CK(_06569_ ), .Q(\ea_wdata[31] ), .QN(_06888_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_1 ( .D(_00270_ ), .CK(_06569_ ), .Q(\ea_wdata[30] ), .QN(_06887_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_10 ( .D(_00271_ ), .CK(_06569_ ), .Q(\ea_wdata[21] ), .QN(_06886_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_11 ( .D(_00272_ ), .CK(_06569_ ), .Q(\ea_wdata[20] ), .QN(_06885_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_12 ( .D(_00273_ ), .CK(_06569_ ), .Q(\ea_wdata[19] ), .QN(_06884_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_13 ( .D(_00274_ ), .CK(_06569_ ), .Q(\ea_wdata[18] ), .QN(_06883_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_14 ( .D(_00275_ ), .CK(_06569_ ), .Q(\ea_wdata[17] ), .QN(_06882_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_15 ( .D(_00276_ ), .CK(_06569_ ), .Q(\ea_wdata[16] ), .QN(_06881_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_16 ( .D(_00277_ ), .CK(_06569_ ), .Q(\ea_wdata[15] ), .QN(_06880_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_17 ( .D(_00278_ ), .CK(_06569_ ), .Q(\ea_wdata[14] ), .QN(_06879_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_18 ( .D(_00279_ ), .CK(_06569_ ), .Q(\ea_wdata[13] ), .QN(_06878_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_19 ( .D(_00280_ ), .CK(_06569_ ), .Q(\ea_wdata[12] ), .QN(_06877_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_2 ( .D(_00281_ ), .CK(_06569_ ), .Q(\ea_wdata[29] ), .QN(_06876_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_20 ( .D(_00282_ ), .CK(_06569_ ), .Q(\ea_wdata[11] ), .QN(_06875_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_21 ( .D(_00283_ ), .CK(_06569_ ), .Q(\ea_wdata[10] ), .QN(_06874_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_22 ( .D(_00284_ ), .CK(_06569_ ), .Q(\ea_wdata[9] ), .QN(_06873_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_23 ( .D(_00285_ ), .CK(_06569_ ), .Q(\ea_wdata[8] ), .QN(_06872_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_24 ( .D(_00286_ ), .CK(_06569_ ), .Q(\ea_wdata[7] ), .QN(_06871_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_25 ( .D(_00287_ ), .CK(_06569_ ), .Q(\ea_wdata[6] ), .QN(_06870_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_26 ( .D(_00288_ ), .CK(_06569_ ), .Q(\ea_wdata[5] ), .QN(_06869_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_27 ( .D(_00289_ ), .CK(_06569_ ), .Q(\ea_wdata[4] ), .QN(_06868_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_28 ( .D(_00290_ ), .CK(_06569_ ), .Q(\ea_wdata[3] ), .QN(_06867_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_29 ( .D(_00291_ ), .CK(_06569_ ), .Q(\ea_wdata[2] ), .QN(_06866_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_3 ( .D(_00292_ ), .CK(_06569_ ), .Q(\ea_wdata[28] ), .QN(_06865_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_30 ( .D(_00293_ ), .CK(_06569_ ), .Q(\ea_wdata[1] ), .QN(_06864_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_31 ( .D(_00294_ ), .CK(_06569_ ), .Q(\ea_wdata[0] ), .QN(_06863_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_4 ( .D(_00295_ ), .CK(_06569_ ), .Q(\ea_wdata[27] ), .QN(_06862_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_5 ( .D(_00296_ ), .CK(_06569_ ), .Q(\ea_wdata[26] ), .QN(_06861_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_6 ( .D(_00297_ ), .CK(_06569_ ), .Q(\ea_wdata[25] ), .QN(_06860_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_7 ( .D(_00298_ ), .CK(_06569_ ), .Q(\ea_wdata[24] ), .QN(_06859_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_8 ( .D(_00299_ ), .CK(_06569_ ), .Q(\ea_wdata[23] ), .QN(_06858_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_9 ( .D(_00300_ ), .CK(_06569_ ), .Q(\ea_wdata[22] ), .QN(_06857_ ) );
DFF_X1 \u_exu.exe_end_$_SDFFE_PP0P__Q ( .D(_00301_ ), .CK(_06567_ ), .Q(exu_valid ), .QN(_06856_ ) );
DFF_X1 \u_exu.exe_start_$_SDFFE_PP0P__Q ( .D(_00302_ ), .CK(_06566_ ), .Q(\u_exu.exe_start ), .QN(_06855_ ) );
DFF_X1 \u_exu.jmpc_ok_$_SDFF_PP0__Q ( .D(_00304_ ), .CK(clock ), .Q(\u_exu.jmpc_ok ), .QN(_06853_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q ( .D(_00303_ ), .CK(_06569_ ), .Q(\ea_addr[31] ), .QN(_06854_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_1 ( .D(_00305_ ), .CK(_06569_ ), .Q(\ea_addr[30] ), .QN(_06852_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_10 ( .D(_00306_ ), .CK(_06569_ ), .Q(\ea_addr[21] ), .QN(_06851_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_11 ( .D(_00307_ ), .CK(_06569_ ), .Q(\ea_addr[20] ), .QN(_06850_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_12 ( .D(_00308_ ), .CK(_06569_ ), .Q(\ea_addr[19] ), .QN(_06849_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_13 ( .D(_00309_ ), .CK(_06569_ ), .Q(\ea_addr[18] ), .QN(_06848_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_14 ( .D(_00310_ ), .CK(_06569_ ), .Q(\ea_addr[17] ), .QN(_06847_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_15 ( .D(_00311_ ), .CK(_06569_ ), .Q(\ea_addr[16] ), .QN(_06846_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_16 ( .D(_00312_ ), .CK(_06569_ ), .Q(\ea_addr[15] ), .QN(_06845_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_17 ( .D(_00313_ ), .CK(_06569_ ), .Q(\ea_addr[14] ), .QN(_06844_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_18 ( .D(_00314_ ), .CK(_06569_ ), .Q(\ea_addr[13] ), .QN(_06843_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_19 ( .D(_00315_ ), .CK(_06569_ ), .Q(\ea_addr[12] ), .QN(_06842_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_2 ( .D(_00316_ ), .CK(_06569_ ), .Q(\ea_addr[29] ), .QN(_06841_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_20 ( .D(_00317_ ), .CK(_06569_ ), .Q(\ea_addr[11] ), .QN(_06840_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_21 ( .D(_00318_ ), .CK(_06569_ ), .Q(\ea_addr[10] ), .QN(_06839_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_22 ( .D(_00319_ ), .CK(_06569_ ), .Q(\ea_addr[9] ), .QN(_06838_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_23 ( .D(_00320_ ), .CK(_06569_ ), .Q(\ea_addr[8] ), .QN(_06837_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_24 ( .D(_00321_ ), .CK(_06569_ ), .Q(\ea_addr[7] ), .QN(_06836_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_25 ( .D(_00322_ ), .CK(_06569_ ), .Q(\ea_addr[6] ), .QN(_06835_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_26 ( .D(_00323_ ), .CK(_06569_ ), .Q(\ea_addr[5] ), .QN(_06834_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_27 ( .D(_00324_ ), .CK(_06569_ ), .Q(\ea_addr[4] ), .QN(_06833_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_28 ( .D(_00325_ ), .CK(_06569_ ), .Q(\ea_addr[3] ), .QN(_06832_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_29 ( .D(_00326_ ), .CK(_06569_ ), .Q(\ea_addr[2] ), .QN(_06831_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_3 ( .D(_00327_ ), .CK(_06569_ ), .Q(\ea_addr[28] ), .QN(_06830_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_30 ( .D(_00328_ ), .CK(_06569_ ), .Q(\ea_addr[1] ), .QN(_06829_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_31 ( .D(_00329_ ), .CK(_06569_ ), .Q(\ea_addr[0] ), .QN(_06828_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_4 ( .D(_00330_ ), .CK(_06569_ ), .Q(\ea_addr[27] ), .QN(_06827_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_5 ( .D(_00331_ ), .CK(_06569_ ), .Q(\ea_addr[26] ), .QN(_06826_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_6 ( .D(_00332_ ), .CK(_06569_ ), .Q(\ea_addr[25] ), .QN(_06825_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_7 ( .D(_00333_ ), .CK(_06569_ ), .Q(\ea_addr[24] ), .QN(_06824_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_8 ( .D(_00334_ ), .CK(_06569_ ), .Q(\ea_addr[23] ), .QN(_06823_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_9 ( .D(_00335_ ), .CK(_06569_ ), .Q(\ea_addr[22] ), .QN(_06822_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q ( .D(_00337_ ), .CK(clock ), .Q(\u_exu.rlock[15] ), .QN(_06820_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_1 ( .D(_00338_ ), .CK(clock ), .Q(\u_exu.rlock[14] ), .QN(_06819_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_10 ( .D(_00339_ ), .CK(clock ), .Q(\u_exu.rlock[5] ), .QN(_06818_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_11 ( .D(_00340_ ), .CK(clock ), .Q(\u_exu.rlock[4] ), .QN(_06817_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_12 ( .D(_00341_ ), .CK(clock ), .Q(\u_exu.rlock[3] ), .QN(_06816_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_13 ( .D(_00342_ ), .CK(clock ), .Q(\u_exu.rlock[2] ), .QN(_06815_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_14 ( .D(_00343_ ), .CK(clock ), .Q(\u_exu.rlock[1] ), .QN(_06814_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_15 ( .D(_00344_ ), .CK(clock ), .Q(\u_exu.rlock[0] ), .QN(_06813_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_2 ( .D(_00345_ ), .CK(clock ), .Q(\u_exu.rlock[13] ), .QN(_06812_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_3 ( .D(_00346_ ), .CK(clock ), .Q(\u_exu.rlock[12] ), .QN(_06811_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_4 ( .D(_00347_ ), .CK(clock ), .Q(\u_exu.rlock[11] ), .QN(_06810_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_5 ( .D(_00348_ ), .CK(clock ), .Q(\u_exu.rlock[10] ), .QN(_06809_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_6 ( .D(_00349_ ), .CK(clock ), .Q(\u_exu.rlock[9] ), .QN(_06808_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_7 ( .D(_00350_ ), .CK(clock ), .Q(\u_exu.rlock[8] ), .QN(_06807_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_8 ( .D(_00351_ ), .CK(clock ), .Q(\u_exu.rlock[7] ), .QN(_06806_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_9 ( .D(_00352_ ), .CK(clock ), .Q(\u_exu.rlock[6] ), .QN(_06805_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q ( .D(_00336_ ), .CK(_06565_ ), .Q(\ca_addr[31] ), .QN(_06821_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_1 ( .D(_00353_ ), .CK(_06565_ ), .Q(\ca_addr[30] ), .QN(_06804_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_10 ( .D(_00354_ ), .CK(_06565_ ), .Q(\ca_addr[21] ), .QN(_06803_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_11 ( .D(_00355_ ), .CK(_06565_ ), .Q(\ca_addr[20] ), .QN(_06802_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_12 ( .D(_00356_ ), .CK(_06565_ ), .Q(\ca_addr[19] ), .QN(_06801_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_13 ( .D(_00357_ ), .CK(_06565_ ), .Q(\ca_addr[18] ), .QN(_06800_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_14 ( .D(_00358_ ), .CK(_06565_ ), .Q(\ca_addr[17] ), .QN(_06799_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_15 ( .D(_00359_ ), .CK(_06565_ ), .Q(\ca_addr[16] ), .QN(_06798_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_16 ( .D(_00360_ ), .CK(_06565_ ), .Q(\ca_addr[15] ), .QN(_06797_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_17 ( .D(_00361_ ), .CK(_06565_ ), .Q(\ca_addr[14] ), .QN(_06796_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_18 ( .D(_00362_ ), .CK(_06565_ ), .Q(\ca_addr[13] ), .QN(_06795_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_19 ( .D(_00363_ ), .CK(_06565_ ), .Q(\ca_addr[12] ), .QN(_06794_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_2 ( .D(_00364_ ), .CK(_06565_ ), .Q(\ca_addr[29] ), .QN(_06793_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_20 ( .D(_00365_ ), .CK(_06565_ ), .Q(\ca_addr[11] ), .QN(_06792_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_21 ( .D(_00366_ ), .CK(_06565_ ), .Q(\ca_addr[10] ), .QN(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_A ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_22 ( .D(_00367_ ), .CK(_06565_ ), .Q(\ca_addr[9] ), .QN(_06791_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_23 ( .D(_00368_ ), .CK(_06565_ ), .Q(\ca_addr[8] ), .QN(io_master_rready_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_24 ( .D(_00369_ ), .CK(_06565_ ), .Q(\ca_addr[7] ), .QN(_06790_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_25 ( .D(_00370_ ), .CK(_06565_ ), .Q(\ca_addr[6] ), .QN(io_master_araddr_$_NOT__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_26 ( .D(_00371_ ), .CK(_06565_ ), .Q(\ca_addr[5] ), .QN(_06789_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_27 ( .D(_00372_ ), .CK(_06565_ ), .Q(\ca_addr[4] ), .QN(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_A ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_3 ( .D(_00373_ ), .CK(_06565_ ), .Q(\ca_addr[28] ), .QN(_06788_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_4 ( .D(_00374_ ), .CK(_06565_ ), .Q(\ca_addr[27] ), .QN(_06787_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_5 ( .D(_00375_ ), .CK(_06565_ ), .Q(\ca_addr[26] ), .QN(_06786_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_6 ( .D(_00376_ ), .CK(_06565_ ), .Q(\ca_addr[25] ), .QN(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_A ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_7 ( .D(_00377_ ), .CK(_06565_ ), .Q(\ca_addr[24] ), .QN(_06785_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_8 ( .D(_00378_ ), .CK(_06565_ ), .Q(\ca_addr[23] ), .QN(_06784_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_9 ( .D(_00379_ ), .CK(_06565_ ), .Q(\ca_addr[22] ), .QN(_07230_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][31] ), .QN(_07231_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][30] ), .QN(_07232_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][21] ), .QN(_07233_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][20] ), .QN(_07234_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][19] ), .QN(_07235_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][18] ), .QN(_07236_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][17] ), .QN(_07237_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][16] ), .QN(_07238_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][15] ), .QN(_07239_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][14] ), .QN(_07240_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][13] ), .QN(_07241_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][12] ), .QN(_07242_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][29] ), .QN(_07243_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][11] ), .QN(_07244_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][10] ), .QN(_07245_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][9] ), .QN(_07246_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][8] ), .QN(_07247_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][7] ), .QN(_07248_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][6] ), .QN(_07249_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][5] ), .QN(_07250_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][4] ), .QN(_07251_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][3] ), .QN(_07252_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][2] ), .QN(_07253_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][28] ), .QN(_07254_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][1] ), .QN(_07255_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][0] ), .QN(_07256_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][27] ), .QN(_07257_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][26] ), .QN(_07258_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][25] ), .QN(_07259_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][24] ), .QN(_07260_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][23] ), .QN(_07261_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06564_ ), .Q(\u_icache.cblocks[0][22] ), .QN(_07262_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][31] ), .QN(_07263_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][30] ), .QN(_07264_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][21] ), .QN(_07265_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][20] ), .QN(_07266_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][19] ), .QN(_07267_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][18] ), .QN(_07268_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][17] ), .QN(_07269_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][16] ), .QN(_07270_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][15] ), .QN(_07271_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][14] ), .QN(_07272_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][13] ), .QN(_07273_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][12] ), .QN(_07274_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][29] ), .QN(_07275_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][11] ), .QN(_07276_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][10] ), .QN(_07277_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][9] ), .QN(_07278_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][8] ), .QN(_07279_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][7] ), .QN(_07280_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][6] ), .QN(_07281_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][5] ), .QN(_07282_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][4] ), .QN(_07283_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][3] ), .QN(_07284_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][2] ), .QN(_07285_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][28] ), .QN(_07286_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][1] ), .QN(_07287_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][0] ), .QN(_07288_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][27] ), .QN(_07289_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][26] ), .QN(_07290_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][25] ), .QN(_07291_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][24] ), .QN(_07292_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][23] ), .QN(_07293_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06563_ ), .Q(\u_icache.cblocks[1][22] ), .QN(_07294_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][31] ), .QN(_07295_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][30] ), .QN(_07296_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][21] ), .QN(_07297_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][20] ), .QN(_07298_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][19] ), .QN(_07299_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][18] ), .QN(_07300_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][17] ), .QN(_07301_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][16] ), .QN(_07302_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][15] ), .QN(_07303_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][14] ), .QN(_07304_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][13] ), .QN(_07305_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][12] ), .QN(_07306_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][29] ), .QN(_07307_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][11] ), .QN(_07308_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][10] ), .QN(_07309_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][9] ), .QN(_07310_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][8] ), .QN(_07311_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][7] ), .QN(_07312_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][6] ), .QN(_07313_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][5] ), .QN(_07314_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][4] ), .QN(_07315_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][3] ), .QN(_07316_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][2] ), .QN(_07317_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][28] ), .QN(_07318_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][1] ), .QN(_07319_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][0] ), .QN(_07320_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][27] ), .QN(_07321_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][26] ), .QN(_07322_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][25] ), .QN(_07323_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][24] ), .QN(_07324_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][23] ), .QN(_07325_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06562_ ), .Q(\u_icache.cblocks[2][22] ), .QN(_07326_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][31] ), .QN(_07327_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][30] ), .QN(_07328_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][21] ), .QN(_07329_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][20] ), .QN(_07330_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][19] ), .QN(_07331_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][18] ), .QN(_07332_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][17] ), .QN(_07333_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][16] ), .QN(_07334_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][15] ), .QN(_07335_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][14] ), .QN(_07336_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][13] ), .QN(_07337_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][12] ), .QN(_07338_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][29] ), .QN(_07339_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][11] ), .QN(_07340_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][10] ), .QN(_07341_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][9] ), .QN(_07342_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][8] ), .QN(_07343_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][7] ), .QN(_07344_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][6] ), .QN(_07345_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][5] ), .QN(_07346_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][4] ), .QN(_07347_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][3] ), .QN(_07348_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][2] ), .QN(_07349_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][28] ), .QN(_07350_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][1] ), .QN(_07351_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][0] ), .QN(_07352_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][27] ), .QN(_07353_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][26] ), .QN(_07354_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][25] ), .QN(_07355_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][24] ), .QN(_07356_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][23] ), .QN(_07357_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06561_ ), .Q(\u_icache.cblocks[3][22] ), .QN(_07358_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][31] ), .QN(_07359_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][30] ), .QN(_07360_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][21] ), .QN(_07361_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][20] ), .QN(_07362_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][19] ), .QN(_07363_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][18] ), .QN(_07364_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][17] ), .QN(_07365_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][16] ), .QN(_07366_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][15] ), .QN(_07367_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][14] ), .QN(_07368_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][13] ), .QN(_07369_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][12] ), .QN(_07370_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][29] ), .QN(_07371_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][11] ), .QN(_07372_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][10] ), .QN(_07373_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][9] ), .QN(_07374_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][8] ), .QN(_07375_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][7] ), .QN(_07376_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][6] ), .QN(_07377_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][5] ), .QN(_07378_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][4] ), .QN(_07379_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][3] ), .QN(_07380_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][2] ), .QN(_07381_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][28] ), .QN(_07382_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][1] ), .QN(_07383_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][0] ), .QN(_07384_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][27] ), .QN(_07385_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][26] ), .QN(_07386_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][25] ), .QN(_07387_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][24] ), .QN(_07388_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][23] ), .QN(_07389_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06560_ ), .Q(\u_icache.cblocks[4][22] ), .QN(_07390_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][31] ), .QN(_07391_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][30] ), .QN(_07392_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][21] ), .QN(_07393_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][20] ), .QN(_07394_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][19] ), .QN(_07395_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][18] ), .QN(_07396_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][17] ), .QN(_07397_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][16] ), .QN(_07398_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][15] ), .QN(_07399_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][14] ), .QN(_07400_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][13] ), .QN(_07401_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][12] ), .QN(_07402_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][29] ), .QN(_07403_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][11] ), .QN(_07404_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][10] ), .QN(_07405_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][9] ), .QN(_07406_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][8] ), .QN(_07407_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][7] ), .QN(_07408_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][6] ), .QN(_07409_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][5] ), .QN(_07410_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][4] ), .QN(_07411_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][3] ), .QN(_07412_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][2] ), .QN(_07413_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][28] ), .QN(_07414_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][1] ), .QN(_07415_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][0] ), .QN(_07416_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][27] ), .QN(_07417_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][26] ), .QN(_07418_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][25] ), .QN(_07419_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][24] ), .QN(_07420_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][23] ), .QN(_07421_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06559_ ), .Q(\u_icache.cblocks[5][22] ), .QN(_07422_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][31] ), .QN(_07423_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][30] ), .QN(_07424_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][21] ), .QN(_07425_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][20] ), .QN(_07426_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][19] ), .QN(_07427_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][18] ), .QN(_07428_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][17] ), .QN(_07429_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][16] ), .QN(_07430_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][15] ), .QN(_07431_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][14] ), .QN(_07432_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][13] ), .QN(_07433_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][12] ), .QN(_07434_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][29] ), .QN(_07435_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][11] ), .QN(_07436_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][10] ), .QN(_07437_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][9] ), .QN(_07438_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][8] ), .QN(_07439_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][7] ), .QN(_07440_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][6] ), .QN(_07441_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][5] ), .QN(_07442_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][4] ), .QN(_07443_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][3] ), .QN(_07444_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][2] ), .QN(_07445_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][28] ), .QN(_07446_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][1] ), .QN(_07447_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][0] ), .QN(_07448_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][27] ), .QN(_07449_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][26] ), .QN(_07450_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][25] ), .QN(_07451_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][24] ), .QN(_07452_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][23] ), .QN(_07453_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06558_ ), .Q(\u_icache.cblocks[6][22] ), .QN(_07454_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q ( .D(\ac_data[31] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][31] ), .QN(_07455_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_1 ( .D(\ac_data[30] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][30] ), .QN(_07456_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_10 ( .D(\ac_data[21] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][21] ), .QN(_07457_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_11 ( .D(\ac_data[20] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][20] ), .QN(_07458_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_12 ( .D(\ac_data[19] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][19] ), .QN(_07459_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_13 ( .D(\ac_data[18] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][18] ), .QN(_07460_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_14 ( .D(\ac_data[17] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][17] ), .QN(_07461_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_15 ( .D(\ac_data[16] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][16] ), .QN(_07462_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_16 ( .D(\ac_data[15] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][15] ), .QN(_07463_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_17 ( .D(\ac_data[14] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][14] ), .QN(_07464_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_18 ( .D(\ac_data[13] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][13] ), .QN(_07465_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_19 ( .D(\ac_data[12] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][12] ), .QN(_07466_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_2 ( .D(\ac_data[29] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][29] ), .QN(_07467_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_20 ( .D(\ac_data[11] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][11] ), .QN(_07468_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_21 ( .D(\ac_data[10] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][10] ), .QN(_07469_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_22 ( .D(\ac_data[9] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][9] ), .QN(_07470_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_23 ( .D(\ac_data[8] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][8] ), .QN(_07471_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_24 ( .D(\ac_data[7] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][7] ), .QN(_07472_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_25 ( .D(\ac_data[6] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][6] ), .QN(_07473_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_26 ( .D(\ac_data[5] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][5] ), .QN(_07474_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_27 ( .D(\ac_data[4] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][4] ), .QN(_07475_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_28 ( .D(\ac_data[3] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][3] ), .QN(_07476_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_29 ( .D(\ac_data[2] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][2] ), .QN(_07477_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_3 ( .D(\ac_data[28] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][28] ), .QN(_07478_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_30 ( .D(\ac_data[1] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][1] ), .QN(_07479_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_31 ( .D(\ac_data[0] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][0] ), .QN(_07480_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_4 ( .D(\ac_data[27] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][27] ), .QN(_07481_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_5 ( .D(\ac_data[26] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][26] ), .QN(_07482_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_6 ( .D(\ac_data[25] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][25] ), .QN(_07483_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_7 ( .D(\ac_data[24] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][24] ), .QN(_07484_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_8 ( .D(\ac_data[23] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][23] ), .QN(_07485_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_9 ( .D(\ac_data[22] ), .CK(_06557_ ), .Q(\u_icache.cblocks[7][22] ), .QN(_06783_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q ( .D(_00380_ ), .CK(_06556_ ), .Q(\cf_inst[31] ), .QN(_06782_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_1 ( .D(_00381_ ), .CK(_06556_ ), .Q(\cf_inst[30] ), .QN(_06781_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_10 ( .D(_00382_ ), .CK(_06556_ ), .Q(\cf_inst[21] ), .QN(_06780_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_11 ( .D(_00383_ ), .CK(_06556_ ), .Q(\cf_inst[20] ), .QN(_06779_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_12 ( .D(_00384_ ), .CK(_06556_ ), .Q(\cf_inst[19] ), .QN(_06778_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_13 ( .D(_00385_ ), .CK(_06556_ ), .Q(\cf_inst[18] ), .QN(_06777_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_14 ( .D(_00386_ ), .CK(_06556_ ), .Q(\cf_inst[17] ), .QN(_06776_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_15 ( .D(_00387_ ), .CK(_06556_ ), .Q(\cf_inst[16] ), .QN(_06775_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_16 ( .D(_00388_ ), .CK(_06556_ ), .Q(\cf_inst[15] ), .QN(_06774_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_17 ( .D(_00389_ ), .CK(_06556_ ), .Q(\cf_inst[14] ), .QN(_06773_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_18 ( .D(_00390_ ), .CK(_06556_ ), .Q(\cf_inst[13] ), .QN(_06772_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_19 ( .D(_00391_ ), .CK(_06556_ ), .Q(\cf_inst[12] ), .QN(_06771_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_2 ( .D(_00392_ ), .CK(_06556_ ), .Q(\cf_inst[29] ), .QN(_06770_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_20 ( .D(_00393_ ), .CK(_06556_ ), .Q(\cf_inst[11] ), .QN(_06769_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_21 ( .D(_00394_ ), .CK(_06556_ ), .Q(\cf_inst[10] ), .QN(_06768_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_22 ( .D(_00395_ ), .CK(_06556_ ), .Q(\cf_inst[9] ), .QN(_06767_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_23 ( .D(_00396_ ), .CK(_06556_ ), .Q(\cf_inst[8] ), .QN(_06766_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_24 ( .D(_00397_ ), .CK(_06556_ ), .Q(\cf_inst[7] ), .QN(_06765_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_25 ( .D(_00398_ ), .CK(_06556_ ), .Q(\cf_inst[6] ), .QN(_06764_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_26 ( .D(_00399_ ), .CK(_06556_ ), .Q(\cf_inst[5] ), .QN(_06763_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_27 ( .D(_00400_ ), .CK(_06556_ ), .Q(\cf_inst[4] ), .QN(_06762_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_28 ( .D(_00401_ ), .CK(_06556_ ), .Q(\cf_inst[3] ), .QN(_06761_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_29 ( .D(_00402_ ), .CK(_06556_ ), .Q(\cf_inst[2] ), .QN(_06760_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_3 ( .D(_00403_ ), .CK(_06556_ ), .Q(\cf_inst[28] ), .QN(_06759_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_30 ( .D(_00404_ ), .CK(_06556_ ), .Q(\cf_inst[1] ), .QN(_06758_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_31 ( .D(_00405_ ), .CK(_06556_ ), .Q(\cf_inst[0] ), .QN(_06757_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_4 ( .D(_00406_ ), .CK(_06556_ ), .Q(\cf_inst[27] ), .QN(_06756_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_5 ( .D(_00407_ ), .CK(_06556_ ), .Q(\cf_inst[26] ), .QN(_06755_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_6 ( .D(_00408_ ), .CK(_06556_ ), .Q(\cf_inst[25] ), .QN(_06754_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_7 ( .D(_00409_ ), .CK(_06556_ ), .Q(\cf_inst[24] ), .QN(_06753_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_8 ( .D(_00410_ ), .CK(_06556_ ), .Q(\cf_inst[23] ), .QN(_06752_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_9 ( .D(_00411_ ), .CK(_06556_ ), .Q(\cf_inst[22] ), .QN(_06751_ ) );
DFF_X1 \u_icache.chvalid_$_SDFFE_PP0P__Q ( .D(_00412_ ), .CK(_06555_ ), .Q(icah_valid ), .QN(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ) );
DFF_X1 \u_icache.count_$_SDFFE_PP0P__Q ( .D(_00413_ ), .CK(_06554_ ), .Q(\u_icache.count[2] ), .QN(_06750_ ) );
DFF_X1 \u_icache.count_$_SDFFE_PP0P__Q_1 ( .D(_00414_ ), .CK(_06554_ ), .Q(\u_icache.count[1] ), .QN(_06749_ ) );
DFF_X1 \u_icache.count_$_SDFFE_PP0P__Q_2 ( .D(_00415_ ), .CK(_06554_ ), .Q(\u_icache.count[0] ), .QN(\u_icache.count_$_NOT__A_Y ) );
DFF_X1 \u_icache.cready_$_SDFF_PP0__Q ( .D(_00416_ ), .CK(clock ), .Q(ifu_ready ), .QN(_07486_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q ( .D(\fc_addr[31] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][26] ), .QN(_06748_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_1 ( .D(\fc_addr[30] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][25] ), .QN(_07487_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_10 ( .D(\fc_addr[21] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][16] ), .QN(_07488_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_11 ( .D(\fc_addr[20] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][15] ), .QN(_07489_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_12 ( .D(\fc_addr[19] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][14] ), .QN(_07490_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_13 ( .D(\fc_addr[18] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][13] ), .QN(_07491_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_14 ( .D(\fc_addr[17] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][12] ), .QN(_07492_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_15 ( .D(\fc_addr[16] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][11] ), .QN(_07493_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_16 ( .D(\fc_addr[15] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][10] ), .QN(_07494_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_17 ( .D(\fc_addr[14] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][9] ), .QN(_07495_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_18 ( .D(\fc_addr[13] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][8] ), .QN(_07496_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_19 ( .D(\fc_addr[12] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][7] ), .QN(_07497_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_2 ( .D(\fc_addr[29] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][24] ), .QN(_07498_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_20 ( .D(\fc_addr[11] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][6] ), .QN(_07499_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_21 ( .D(\fc_addr[10] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][5] ), .QN(_07500_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_22 ( .D(\fc_addr[9] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][4] ), .QN(_07501_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_23 ( .D(\fc_addr[8] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][3] ), .QN(_07502_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_24 ( .D(\fc_addr[7] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][2] ), .QN(_07503_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_25 ( .D(\fc_addr[6] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][1] ), .QN(_07504_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_26 ( .D(\fc_addr[5] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][0] ), .QN(_07505_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_3 ( .D(\fc_addr[28] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][23] ), .QN(_07506_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_4 ( .D(\fc_addr[27] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][22] ), .QN(_07507_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_5 ( .D(\fc_addr[26] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][21] ), .QN(_07508_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_6 ( .D(\fc_addr[25] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][20] ), .QN(_07509_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_7 ( .D(\fc_addr[24] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][19] ), .QN(_07510_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_8 ( .D(\fc_addr[23] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][18] ), .QN(_07511_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_9 ( .D(\fc_addr[22] ), .CK(_06553_ ), .Q(\u_icache.ctags[0][17] ), .QN(_07512_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q ( .D(\fc_addr[31] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][26] ), .QN(_07513_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_1 ( .D(\fc_addr[30] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][25] ), .QN(_07514_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_10 ( .D(\fc_addr[21] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][16] ), .QN(_07515_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_11 ( .D(\fc_addr[20] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][15] ), .QN(_07516_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_12 ( .D(\fc_addr[19] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][14] ), .QN(_07517_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_13 ( .D(\fc_addr[18] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][13] ), .QN(_07518_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_14 ( .D(\fc_addr[17] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][12] ), .QN(_07519_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_15 ( .D(\fc_addr[16] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][11] ), .QN(_07520_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_16 ( .D(\fc_addr[15] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][10] ), .QN(_07521_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_17 ( .D(\fc_addr[14] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][9] ), .QN(_07522_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_18 ( .D(\fc_addr[13] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][8] ), .QN(_07523_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_19 ( .D(\fc_addr[12] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][7] ), .QN(_07524_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_2 ( .D(\fc_addr[29] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][24] ), .QN(_07525_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_20 ( .D(\fc_addr[11] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][6] ), .QN(_07526_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_21 ( .D(\fc_addr[10] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][5] ), .QN(_07527_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_22 ( .D(\fc_addr[9] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][4] ), .QN(_07528_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_23 ( .D(\fc_addr[8] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][3] ), .QN(_07529_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_24 ( .D(\fc_addr[7] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][2] ), .QN(_07530_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_25 ( .D(\fc_addr[6] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][1] ), .QN(_07531_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_26 ( .D(\fc_addr[5] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][0] ), .QN(_07532_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_3 ( .D(\fc_addr[28] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][23] ), .QN(_07533_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_4 ( .D(\fc_addr[27] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][22] ), .QN(_07534_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_5 ( .D(\fc_addr[26] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][21] ), .QN(_07535_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_6 ( .D(\fc_addr[25] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][20] ), .QN(_07536_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_7 ( .D(\fc_addr[24] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][19] ), .QN(_07537_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_8 ( .D(\fc_addr[23] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][18] ), .QN(_07538_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_9 ( .D(\fc_addr[22] ), .CK(_06552_ ), .Q(\u_icache.ctags[1][17] ), .QN(_06747_ ) );
DFF_X1 \u_icache.cvalids_$_SDFFE_PP0P__Q ( .D(_00417_ ), .CK(_06551_ ), .Q(\u_icache.cvalids[1] ), .QN(_06746_ ) );
DFF_X1 \u_icache.cvalids_$_SDFFE_PP0P__Q_1 ( .D(_00418_ ), .CK(_06551_ ), .Q(\u_icache.cvalids[0] ), .QN(_06745_ ) );
DFF_X1 \u_icache.ended_$_SDFFE_PP0P__Q ( .D(_00419_ ), .CK(_06550_ ), .Q(\u_icache.ended ), .QN(_06744_ ) );
DFF_X1 \u_idu.decode_ok_$_SDFFE_PP0P__Q ( .D(_00420_ ), .CK(_06549_ ), .Q(exe_valid ), .QN(_06743_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q ( .D(_00421_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[31] ), .QN(_06742_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_1 ( .D(_00422_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[30] ), .QN(\u_exu.opt_$_NOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_10 ( .D(_00423_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[21] ), .QN(_06741_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_11 ( .D(_00424_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[20] ), .QN(\u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_12 ( .D(_00425_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[19] ), .QN(_06740_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_13 ( .D(_00426_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[18] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_14 ( .D(_00427_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[17] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_1_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_15 ( .D(_00428_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[16] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_16 ( .D(_00429_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[15] ), .QN(_06739_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_17 ( .D(_00430_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[14] ), .QN(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_18 ( .D(_00431_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[13] ), .QN(de_ard_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_19 ( .D(_00432_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[12] ), .QN(_06738_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_2 ( .D(_00433_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[29] ), .QN(_06737_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_20 ( .D(_00434_ ), .CK(_06548_ ), .Q(\u_idu.imm_branch[4] ), .QN(_06736_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_21 ( .D(_00435_ ), .CK(_06548_ ), .Q(\u_idu.imm_branch[3] ), .QN(_06735_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_22 ( .D(_00436_ ), .CK(_06548_ ), .Q(\u_idu.imm_branch[2] ), .QN(_06734_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_23 ( .D(_00437_ ), .CK(_06548_ ), .Q(\u_idu.imm_branch[1] ), .QN(_06733_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_24 ( .D(_00438_ ), .CK(_06548_ ), .Q(\u_idu.imm_branch[11] ), .QN(_06732_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_25 ( .D(_00439_ ), .CK(_06548_ ), .Q(\u_idu.inst[6] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_26 ( .D(_00440_ ), .CK(_06548_ ), .Q(\u_idu.inst[5] ), .QN(_06731_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_27 ( .D(_00441_ ), .CK(_06548_ ), .Q(\u_idu.inst[4] ), .QN(_06730_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_28 ( .D(_00442_ ), .CK(_06548_ ), .Q(\u_idu.inst[3] ), .QN(_06729_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_29 ( .D(_00443_ ), .CK(_06548_ ), .Q(\u_idu.inst[2] ), .QN(_06728_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_3 ( .D(_00444_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[28] ), .QN(_06727_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_30 ( .D(_00445_ ), .CK(_06548_ ), .Q(\u_idu.inst[1] ), .QN(_06726_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_31 ( .D(_00446_ ), .CK(_06548_ ), .Q(\u_idu.inst[0] ), .QN(_06725_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_4 ( .D(_00447_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[27] ), .QN(_06724_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_5 ( .D(_00448_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[26] ), .QN(_06723_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_6 ( .D(_00449_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[25] ), .QN(_06722_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_7 ( .D(_00450_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[24] ), .QN(_06721_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_8 ( .D(_00451_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[23] ), .QN(_06720_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_9 ( .D(_00452_ ), .CK(_06548_ ), .Q(\u_idu.imm_auipc_lui[22] ), .QN(_06719_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q ( .D(_00453_ ), .CK(_06548_ ), .Q(\de_pc[31] ), .QN(_06718_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00454_ ), .CK(_06548_ ), .Q(\de_pc[30] ), .QN(_06717_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00455_ ), .CK(_06548_ ), .Q(\de_pc[21] ), .QN(_06716_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00456_ ), .CK(_06548_ ), .Q(\de_pc[20] ), .QN(_06715_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00457_ ), .CK(_06548_ ), .Q(\de_pc[19] ), .QN(_06714_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00458_ ), .CK(_06548_ ), .Q(\de_pc[18] ), .QN(_06713_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00459_ ), .CK(_06548_ ), .Q(\de_pc[17] ), .QN(_06712_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00460_ ), .CK(_06548_ ), .Q(\de_pc[16] ), .QN(_06711_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00461_ ), .CK(_06548_ ), .Q(\de_pc[15] ), .QN(_06710_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00462_ ), .CK(_06548_ ), .Q(\de_pc[14] ), .QN(_06709_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00463_ ), .CK(_06548_ ), .Q(\de_pc[13] ), .QN(_06708_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00464_ ), .CK(_06548_ ), .Q(\de_pc[12] ), .QN(_06707_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00465_ ), .CK(_06548_ ), .Q(\de_pc[29] ), .QN(_06706_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00466_ ), .CK(_06548_ ), .Q(\de_pc[11] ), .QN(_06705_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00467_ ), .CK(_06548_ ), .Q(\de_pc[10] ), .QN(_06704_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00468_ ), .CK(_06548_ ), .Q(\de_pc[9] ), .QN(_06703_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00469_ ), .CK(_06548_ ), .Q(\de_pc[8] ), .QN(_06702_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00470_ ), .CK(_06548_ ), .Q(\de_pc[7] ), .QN(_06701_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00471_ ), .CK(_06548_ ), .Q(\de_pc[6] ), .QN(_06700_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00472_ ), .CK(_06548_ ), .Q(\de_pc[5] ), .QN(_06699_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00473_ ), .CK(_06548_ ), .Q(\de_pc[4] ), .QN(_06698_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00474_ ), .CK(_06548_ ), .Q(\de_pc[3] ), .QN(_06697_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00475_ ), .CK(_06548_ ), .Q(\de_pc[2] ), .QN(_06696_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00476_ ), .CK(_06548_ ), .Q(\de_pc[28] ), .QN(_06695_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00477_ ), .CK(_06548_ ), .Q(\de_pc[1] ), .QN(_06694_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_31 ( .D(_00478_ ), .CK(_06548_ ), .Q(\de_pc[0] ), .QN(_06693_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00479_ ), .CK(_06548_ ), .Q(\de_pc[27] ), .QN(_06692_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00480_ ), .CK(_06548_ ), .Q(\de_pc[26] ), .QN(_06691_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00481_ ), .CK(_06548_ ), .Q(\de_pc[25] ), .QN(_06690_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00482_ ), .CK(_06548_ ), .Q(\de_pc[24] ), .QN(_06689_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00483_ ), .CK(_06548_ ), .Q(\de_pc[23] ), .QN(_06688_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00484_ ), .CK(_06548_ ), .Q(\de_pc[22] ), .QN(_06687_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q ( .D(_00485_ ), .CK(_06547_ ), .Q(\fd_inst[31] ), .QN(_06686_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_1 ( .D(_00486_ ), .CK(_06547_ ), .Q(\fd_inst[30] ), .QN(_06685_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_10 ( .D(_00487_ ), .CK(_06547_ ), .Q(\fd_inst[21] ), .QN(_06684_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_11 ( .D(_00488_ ), .CK(_06547_ ), .Q(\fd_inst[20] ), .QN(_06683_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_12 ( .D(_00489_ ), .CK(_06547_ ), .Q(\fd_inst[19] ), .QN(_06682_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_13 ( .D(_00490_ ), .CK(_06547_ ), .Q(\fd_inst[18] ), .QN(_06681_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_14 ( .D(_00491_ ), .CK(_06547_ ), .Q(\fd_inst[17] ), .QN(_06680_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_15 ( .D(_00492_ ), .CK(_06547_ ), .Q(\fd_inst[16] ), .QN(_06679_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_16 ( .D(_00493_ ), .CK(_06547_ ), .Q(\fd_inst[15] ), .QN(_06678_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_17 ( .D(_00494_ ), .CK(_06547_ ), .Q(\fd_inst[14] ), .QN(_06677_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_18 ( .D(_00495_ ), .CK(_06547_ ), .Q(\fd_inst[13] ), .QN(_06676_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_19 ( .D(_00496_ ), .CK(_06547_ ), .Q(\fd_inst[12] ), .QN(_06675_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_2 ( .D(_00497_ ), .CK(_06547_ ), .Q(\fd_inst[29] ), .QN(_06674_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_20 ( .D(_00498_ ), .CK(_06547_ ), .Q(\fd_inst[11] ), .QN(_06673_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_21 ( .D(_00499_ ), .CK(_06547_ ), .Q(\fd_inst[10] ), .QN(_06672_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_22 ( .D(_00500_ ), .CK(_06547_ ), .Q(\fd_inst[9] ), .QN(_06671_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_23 ( .D(_00501_ ), .CK(_06547_ ), .Q(\fd_inst[8] ), .QN(_06670_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_24 ( .D(_00502_ ), .CK(_06547_ ), .Q(\fd_inst[7] ), .QN(_06669_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_25 ( .D(_00503_ ), .CK(_06547_ ), .Q(\fd_inst[6] ), .QN(_06668_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_26 ( .D(_00504_ ), .CK(_06547_ ), .Q(\fd_inst[5] ), .QN(_06667_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_27 ( .D(_00505_ ), .CK(_06547_ ), .Q(\fd_inst[4] ), .QN(_06666_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_28 ( .D(_00506_ ), .CK(_06547_ ), .Q(\fd_inst[3] ), .QN(_06665_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_29 ( .D(_00507_ ), .CK(_06547_ ), .Q(\fd_inst[2] ), .QN(_06664_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_3 ( .D(_00508_ ), .CK(_06547_ ), .Q(\fd_inst[28] ), .QN(_06663_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_30 ( .D(_00509_ ), .CK(_06547_ ), .Q(\fd_inst[1] ), .QN(_06662_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_31 ( .D(_00510_ ), .CK(_06547_ ), .Q(\fd_inst[0] ), .QN(_06661_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_4 ( .D(_00511_ ), .CK(_06547_ ), .Q(\fd_inst[27] ), .QN(_06660_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_5 ( .D(_00512_ ), .CK(_06547_ ), .Q(\fd_inst[26] ), .QN(_06659_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_6 ( .D(_00513_ ), .CK(_06547_ ), .Q(\fd_inst[25] ), .QN(_06658_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_7 ( .D(_00514_ ), .CK(_06547_ ), .Q(\fd_inst[24] ), .QN(_06657_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_8 ( .D(_00515_ ), .CK(_06547_ ), .Q(\fd_inst[23] ), .QN(_06656_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_9 ( .D(_00516_ ), .CK(_06547_ ), .Q(\fd_inst[22] ), .QN(_06655_ ) );
DFF_X1 \u_ifu.inst_ok_$_SDFFE_PP0P__Q ( .D(_00517_ ), .CK(_06546_ ), .Q(idu_ready ), .QN(_06654_ ) );
DFF_X1 \u_ifu.jpc_ok_$_SDFFE_PP0P__Q ( .D(_00518_ ), .CK(_06545_ ), .Q(\u_ifu.jpc_ok ), .QN(\u_ifu.jpc_ok_$_NOT__A_Y ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q ( .D(_00519_ ), .CK(_06544_ ), .Q(\fc_addr[30] ), .QN(_06653_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_1 ( .D(_00520_ ), .CK(_06544_ ), .Q(\fc_addr[29] ), .QN(_06652_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_10 ( .D(_00521_ ), .CK(_06544_ ), .Q(\fc_addr[20] ), .QN(_06651_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_11 ( .D(_00522_ ), .CK(_06544_ ), .Q(\fc_addr[19] ), .QN(_06650_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_12 ( .D(_00523_ ), .CK(_06544_ ), .Q(\fc_addr[18] ), .QN(_06649_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_13 ( .D(_00524_ ), .CK(_06544_ ), .Q(\fc_addr[17] ), .QN(_06648_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_14 ( .D(_00525_ ), .CK(_06544_ ), .Q(\fc_addr[16] ), .QN(_06647_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_15 ( .D(_00526_ ), .CK(_06544_ ), .Q(\fc_addr[15] ), .QN(_06646_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_16 ( .D(_00527_ ), .CK(_06544_ ), .Q(\fc_addr[14] ), .QN(_06645_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_17 ( .D(_00528_ ), .CK(_06544_ ), .Q(\fc_addr[13] ), .QN(_06644_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_18 ( .D(_00529_ ), .CK(_06544_ ), .Q(\fc_addr[12] ), .QN(_06643_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_19 ( .D(_00530_ ), .CK(_06544_ ), .Q(\fc_addr[11] ), .QN(_06642_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_2 ( .D(_00531_ ), .CK(_06544_ ), .Q(\fc_addr[28] ), .QN(_06641_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_20 ( .D(_00532_ ), .CK(_06544_ ), .Q(\fc_addr[10] ), .QN(_06640_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_21 ( .D(_00533_ ), .CK(_06544_ ), .Q(\fc_addr[9] ), .QN(_06639_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_22 ( .D(_00534_ ), .CK(_06544_ ), .Q(\fc_addr[8] ), .QN(_06638_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_23 ( .D(_00535_ ), .CK(_06544_ ), .Q(\fc_addr[7] ), .QN(_06637_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_24 ( .D(_00536_ ), .CK(_06544_ ), .Q(\fc_addr[6] ), .QN(_06636_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_25 ( .D(_00537_ ), .CK(_06544_ ), .Q(\fc_addr[5] ), .QN(_06635_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_26 ( .D(_00538_ ), .CK(_06544_ ), .Q(\fc_addr[4] ), .QN(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D ( .D(_00540_ ), .CK(clock ), .Q(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .QN(_06633_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_27 ( .D(_00539_ ), .CK(_06544_ ), .Q(\fc_addr[3] ), .QN(_06634_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_28 ( .D(_00541_ ), .CK(_06544_ ), .Q(\fc_addr[2] ), .QN(\u_ifu.pc_$_SDFFE_PP0N__Q_28_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_3 ( .D(_00542_ ), .CK(_06544_ ), .Q(\fc_addr[27] ), .QN(_06632_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_4 ( .D(_00543_ ), .CK(_06544_ ), .Q(\fc_addr[26] ), .QN(_06631_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_5 ( .D(_00544_ ), .CK(_06544_ ), .Q(\fc_addr[25] ), .QN(_06630_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_6 ( .D(_00545_ ), .CK(_06544_ ), .Q(\fc_addr[24] ), .QN(_06629_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_7 ( .D(_00546_ ), .CK(_06544_ ), .Q(\fc_addr[23] ), .QN(_06628_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_8 ( .D(_00547_ ), .CK(_06544_ ), .Q(\fc_addr[22] ), .QN(_06627_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_9 ( .D(_00548_ ), .CK(_06544_ ), .Q(\fc_addr[21] ), .QN(_06626_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0P__Q ( .D(_00549_ ), .CK(_06543_ ), .Q(\fc_addr[1] ), .QN(_06625_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00550_ ), .CK(_06543_ ), .Q(\fc_addr[0] ), .QN(_06624_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP1N__Q ( .D(_00551_ ), .CK(_06544_ ), .Q(\fc_addr[31] ), .QN(_06623_ ) );
DFF_X1 \u_lsu.arvalid_$_SDFFE_PP0P__Q ( .D(_00552_ ), .CK(_06542_ ), .Q(\u_lsu.arvalid ), .QN(_06622_ ) );
DFF_X1 \u_lsu.awvalid_$_SDFFE_PP0P__Q ( .D(_00553_ ), .CK(_06541_ ), .Q(io_master_awvalid ), .QN(_06621_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q ( .D(_00554_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[7] ), .QN(_06620_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_1 ( .D(_00555_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[6] ), .QN(_06619_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_2 ( .D(_00556_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[5] ), .QN(_06618_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_3 ( .D(_00557_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[4] ), .QN(_06617_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_4 ( .D(_00558_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[3] ), .QN(_06616_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_5 ( .D(_00559_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[2] ), .QN(_06615_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_6 ( .D(_00560_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[1] ), .QN(_06614_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_7 ( .D(_00561_ ), .CK(_06540_ ), .Q(\u_lsu.rcount[0] ), .QN(_06613_ ) );
DFF_X1 \u_lsu.reading_$_SDFFE_PP0P__Q ( .D(_00552_ ), .CK(_06539_ ), .Q(\u_lsu.reading ), .QN(_06612_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q ( .D(_00562_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[63] ), .QN(_06610_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_1 ( .D(_00563_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[62] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_10 ( .D(_00564_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[53] ), .QN(_06609_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_11 ( .D(_00565_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[52] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_10_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_12 ( .D(_00566_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[51] ), .QN(_06608_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_13 ( .D(_00567_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[50] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_14 ( .D(_00568_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[49] ), .QN(_06607_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_15 ( .D(_00569_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[48] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_16 ( .D(_00570_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[47] ), .QN(_06606_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_17 ( .D(_00571_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[46] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_18 ( .D(_00572_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[45] ), .QN(_06605_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_19 ( .D(_00573_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[44] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_18_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_2 ( .D(_00574_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[61] ), .QN(_06604_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_20 ( .D(_00575_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[43] ), .QN(_06603_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_21 ( .D(_00576_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[42] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_22 ( .D(_00577_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[41] ), .QN(_06602_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_23 ( .D(_00578_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[40] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_24 ( .D(_00579_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[39] ), .QN(_06601_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_25 ( .D(_00580_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[38] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_26 ( .D(_00581_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[37] ), .QN(_06600_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_27 ( .D(_00582_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[36] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_26_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_28 ( .D(_00583_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[35] ), .QN(_06599_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_29 ( .D(_00584_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[34] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_28_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_3 ( .D(_00585_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[60] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_30 ( .D(_00586_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[33] ), .QN(_06598_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_31 ( .D(_00587_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[32] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_32 ( .D(_00588_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[31] ), .QN(_06597_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_33 ( .D(_00589_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[30] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_31_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_34 ( .D(_00590_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[29] ), .QN(_06596_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_35 ( .D(_00591_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[28] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_36 ( .D(_00592_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[27] ), .QN(_06595_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_37 ( .D(_00593_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[26] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_38 ( .D(_00594_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[25] ), .QN(_06594_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_39 ( .D(_00595_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[24] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_4 ( .D(_00596_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[59] ), .QN(_06593_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_40 ( .D(_00597_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[23] ), .QN(_06592_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_41 ( .D(_00598_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[22] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_39_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_42 ( .D(_00599_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[21] ), .QN(_06591_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_43 ( .D(_00600_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[20] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_44 ( .D(_00601_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[19] ), .QN(_06590_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_45 ( .D(_00602_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[18] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_46 ( .D(_00603_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[17] ), .QN(_06589_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_47 ( .D(_00604_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[16] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_48 ( .D(_00605_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[15] ), .QN(_06588_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_49 ( .D(_00606_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[14] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_5 ( .D(_00607_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[58] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_50 ( .D(_00608_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[13] ), .QN(_06587_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_51 ( .D(_00609_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[12] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_52 ( .D(_00610_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[11] ), .QN(_06586_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_53 ( .D(_00611_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[10] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_54 ( .D(_00612_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[9] ), .QN(_06585_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_55 ( .D(_00613_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[8] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_56 ( .D(_00614_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[7] ), .QN(_06584_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_57 ( .D(_00615_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[6] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_58 ( .D(_00616_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[5] ), .QN(_06583_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_59 ( .D(_00617_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[4] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_6 ( .D(_00618_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[57] ), .QN(_06582_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_60 ( .D(_00619_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[3] ), .QN(_06581_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_61 ( .D(_00620_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[2] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_62 ( .D(_00621_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[1] ), .QN(_06580_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63 ( .D(_00622_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[0] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D[0] ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_7 ( .D(_00623_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[56] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_8 ( .D(_00624_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[55] ), .QN(_06579_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_9 ( .D(_00625_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime[54] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_8_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.tvalid_$_SDFF_PP0__Q ( .D(_00626_ ), .CK(clock ), .Q(\u_lsu.rvalid_clint ), .QN(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \u_lsu.wlast_$_SDFFE_PP0P__Q ( .D(_00553_ ), .CK(_06538_ ), .Q(io_master_wlast ), .QN(_06611_ ) );
DFF_X1 \u_lsu.writing_$_SDFFE_PP0P__Q ( .D(_00553_ ), .CK(_06537_ ), .Q(\u_lsu.writing ), .QN(_07539_ ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06536_ ), .Q(\u_reg.rf[10][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06536_ ), .Q(\u_reg.rf[10][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06536_ ), .Q(\u_reg.rf[10][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06536_ ), .Q(\u_reg.rf[10][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06536_ ), .Q(\u_reg.rf[10][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06536_ ), .Q(\u_reg.rf[10][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06536_ ), .Q(\u_reg.rf[10][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06536_ ), .Q(\u_reg.rf[10][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06536_ ), .Q(\u_reg.rf[10][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06536_ ), .Q(\u_reg.rf[10][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06536_ ), .Q(\u_reg.rf[10][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06536_ ), .Q(\u_reg.rf[10][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06536_ ), .Q(\u_reg.rf[10][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06536_ ), .Q(\u_reg.rf[10][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06536_ ), .Q(\u_reg.rf[10][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06536_ ), .Q(\u_reg.rf[10][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06536_ ), .Q(\u_reg.rf[10][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06536_ ), .Q(\u_reg.rf[10][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06536_ ), .Q(\u_reg.rf[10][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06536_ ), .Q(\u_reg.rf[10][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06536_ ), .Q(\u_reg.rf[10][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06536_ ), .Q(\u_reg.rf[10][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06536_ ), .Q(\u_reg.rf[10][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06536_ ), .Q(\u_reg.rf[10][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06536_ ), .Q(\u_reg.rf[10][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06536_ ), .Q(\u_reg.rf[10][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06536_ ), .Q(\u_reg.rf[10][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06536_ ), .Q(\u_reg.rf[10][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06536_ ), .Q(\u_reg.rf[10][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06536_ ), .Q(\u_reg.rf[10][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06536_ ), .Q(\u_reg.rf[10][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06536_ ), .Q(\u_reg.rf[10][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06535_ ), .Q(\u_reg.rf[11][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06535_ ), .Q(\u_reg.rf[11][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06535_ ), .Q(\u_reg.rf[11][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06535_ ), .Q(\u_reg.rf[11][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06535_ ), .Q(\u_reg.rf[11][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06535_ ), .Q(\u_reg.rf[11][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06535_ ), .Q(\u_reg.rf[11][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06535_ ), .Q(\u_reg.rf[11][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06535_ ), .Q(\u_reg.rf[11][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06535_ ), .Q(\u_reg.rf[11][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06535_ ), .Q(\u_reg.rf[11][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06535_ ), .Q(\u_reg.rf[11][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06535_ ), .Q(\u_reg.rf[11][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06535_ ), .Q(\u_reg.rf[11][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06535_ ), .Q(\u_reg.rf[11][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06535_ ), .Q(\u_reg.rf[11][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06535_ ), .Q(\u_reg.rf[11][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06535_ ), .Q(\u_reg.rf[11][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06535_ ), .Q(\u_reg.rf[11][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06535_ ), .Q(\u_reg.rf[11][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06535_ ), .Q(\u_reg.rf[11][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06535_ ), .Q(\u_reg.rf[11][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06535_ ), .Q(\u_reg.rf[11][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06535_ ), .Q(\u_reg.rf[11][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06535_ ), .Q(\u_reg.rf[11][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06535_ ), .Q(\u_reg.rf[11][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06535_ ), .Q(\u_reg.rf[11][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06535_ ), .Q(\u_reg.rf[11][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06535_ ), .Q(\u_reg.rf[11][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06535_ ), .Q(\u_reg.rf[11][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06535_ ), .Q(\u_reg.rf[11][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06535_ ), .Q(\u_reg.rf[11][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06534_ ), .Q(\u_reg.rf[12][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06534_ ), .Q(\u_reg.rf[12][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06534_ ), .Q(\u_reg.rf[12][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06534_ ), .Q(\u_reg.rf[12][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06534_ ), .Q(\u_reg.rf[12][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06534_ ), .Q(\u_reg.rf[12][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06534_ ), .Q(\u_reg.rf[12][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06534_ ), .Q(\u_reg.rf[12][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06534_ ), .Q(\u_reg.rf[12][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06534_ ), .Q(\u_reg.rf[12][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06534_ ), .Q(\u_reg.rf[12][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06534_ ), .Q(\u_reg.rf[12][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06534_ ), .Q(\u_reg.rf[12][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06534_ ), .Q(\u_reg.rf[12][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06534_ ), .Q(\u_reg.rf[12][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06534_ ), .Q(\u_reg.rf[12][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06534_ ), .Q(\u_reg.rf[12][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06534_ ), .Q(\u_reg.rf[12][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06534_ ), .Q(\u_reg.rf[12][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06534_ ), .Q(\u_reg.rf[12][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06534_ ), .Q(\u_reg.rf[12][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06534_ ), .Q(\u_reg.rf[12][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06534_ ), .Q(\u_reg.rf[12][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06534_ ), .Q(\u_reg.rf[12][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06534_ ), .Q(\u_reg.rf[12][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06534_ ), .Q(\u_reg.rf[12][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06534_ ), .Q(\u_reg.rf[12][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06534_ ), .Q(\u_reg.rf[12][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06534_ ), .Q(\u_reg.rf[12][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06534_ ), .Q(\u_reg.rf[12][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06534_ ), .Q(\u_reg.rf[12][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06534_ ), .Q(\u_reg.rf[12][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06533_ ), .Q(\u_reg.rf[13][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06533_ ), .Q(\u_reg.rf[13][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06533_ ), .Q(\u_reg.rf[13][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06533_ ), .Q(\u_reg.rf[13][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06533_ ), .Q(\u_reg.rf[13][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06533_ ), .Q(\u_reg.rf[13][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06533_ ), .Q(\u_reg.rf[13][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06533_ ), .Q(\u_reg.rf[13][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06533_ ), .Q(\u_reg.rf[13][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06533_ ), .Q(\u_reg.rf[13][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06533_ ), .Q(\u_reg.rf[13][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06533_ ), .Q(\u_reg.rf[13][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06533_ ), .Q(\u_reg.rf[13][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06533_ ), .Q(\u_reg.rf[13][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06533_ ), .Q(\u_reg.rf[13][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06533_ ), .Q(\u_reg.rf[13][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06533_ ), .Q(\u_reg.rf[13][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06533_ ), .Q(\u_reg.rf[13][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06533_ ), .Q(\u_reg.rf[13][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06533_ ), .Q(\u_reg.rf[13][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06533_ ), .Q(\u_reg.rf[13][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06533_ ), .Q(\u_reg.rf[13][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06533_ ), .Q(\u_reg.rf[13][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06533_ ), .Q(\u_reg.rf[13][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06533_ ), .Q(\u_reg.rf[13][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06533_ ), .Q(\u_reg.rf[13][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06533_ ), .Q(\u_reg.rf[13][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06533_ ), .Q(\u_reg.rf[13][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06533_ ), .Q(\u_reg.rf[13][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06533_ ), .Q(\u_reg.rf[13][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06533_ ), .Q(\u_reg.rf[13][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06533_ ), .Q(\u_reg.rf[13][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06532_ ), .Q(\u_reg.rf[14][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06532_ ), .Q(\u_reg.rf[14][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06532_ ), .Q(\u_reg.rf[14][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06532_ ), .Q(\u_reg.rf[14][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06532_ ), .Q(\u_reg.rf[14][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06532_ ), .Q(\u_reg.rf[14][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06532_ ), .Q(\u_reg.rf[14][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06532_ ), .Q(\u_reg.rf[14][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06532_ ), .Q(\u_reg.rf[14][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06532_ ), .Q(\u_reg.rf[14][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06532_ ), .Q(\u_reg.rf[14][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06532_ ), .Q(\u_reg.rf[14][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06532_ ), .Q(\u_reg.rf[14][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06532_ ), .Q(\u_reg.rf[14][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06532_ ), .Q(\u_reg.rf[14][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06532_ ), .Q(\u_reg.rf[14][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06532_ ), .Q(\u_reg.rf[14][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06532_ ), .Q(\u_reg.rf[14][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06532_ ), .Q(\u_reg.rf[14][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06532_ ), .Q(\u_reg.rf[14][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06532_ ), .Q(\u_reg.rf[14][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06532_ ), .Q(\u_reg.rf[14][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06532_ ), .Q(\u_reg.rf[14][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06532_ ), .Q(\u_reg.rf[14][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06532_ ), .Q(\u_reg.rf[14][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06532_ ), .Q(\u_reg.rf[14][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06532_ ), .Q(\u_reg.rf[14][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06532_ ), .Q(\u_reg.rf[14][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06532_ ), .Q(\u_reg.rf[14][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06532_ ), .Q(\u_reg.rf[14][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06532_ ), .Q(\u_reg.rf[14][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06532_ ), .Q(\u_reg.rf[14][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06531_ ), .Q(\u_reg.rf[15][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06531_ ), .Q(\u_reg.rf[15][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06531_ ), .Q(\u_reg.rf[15][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06531_ ), .Q(\u_reg.rf[15][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06531_ ), .Q(\u_reg.rf[15][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06531_ ), .Q(\u_reg.rf[15][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06531_ ), .Q(\u_reg.rf[15][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06531_ ), .Q(\u_reg.rf[15][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06531_ ), .Q(\u_reg.rf[15][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06531_ ), .Q(\u_reg.rf[15][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06531_ ), .Q(\u_reg.rf[15][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06531_ ), .Q(\u_reg.rf[15][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06531_ ), .Q(\u_reg.rf[15][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06531_ ), .Q(\u_reg.rf[15][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06531_ ), .Q(\u_reg.rf[15][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06531_ ), .Q(\u_reg.rf[15][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06531_ ), .Q(\u_reg.rf[15][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06531_ ), .Q(\u_reg.rf[15][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06531_ ), .Q(\u_reg.rf[15][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06531_ ), .Q(\u_reg.rf[15][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06531_ ), .Q(\u_reg.rf[15][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06531_ ), .Q(\u_reg.rf[15][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06531_ ), .Q(\u_reg.rf[15][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06531_ ), .Q(\u_reg.rf[15][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06531_ ), .Q(\u_reg.rf[15][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06531_ ), .Q(\u_reg.rf[15][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06531_ ), .Q(\u_reg.rf[15][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06531_ ), .Q(\u_reg.rf[15][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06531_ ), .Q(\u_reg.rf[15][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06531_ ), .Q(\u_reg.rf[15][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06531_ ), .Q(\u_reg.rf[15][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06531_ ), .Q(\u_reg.rf[15][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06530_ ), .Q(\u_reg.rf[1][31] ), .QN(_07540_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06530_ ), .Q(\u_reg.rf[1][30] ), .QN(_07541_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06530_ ), .Q(\u_reg.rf[1][21] ), .QN(_07542_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06530_ ), .Q(\u_reg.rf[1][20] ), .QN(_07543_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06530_ ), .Q(\u_reg.rf[1][19] ), .QN(_07544_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06530_ ), .Q(\u_reg.rf[1][18] ), .QN(_07545_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06530_ ), .Q(\u_reg.rf[1][17] ), .QN(_07546_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06530_ ), .Q(\u_reg.rf[1][16] ), .QN(_07547_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06530_ ), .Q(\u_reg.rf[1][15] ), .QN(_07548_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06530_ ), .Q(\u_reg.rf[1][14] ), .QN(_07549_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06530_ ), .Q(\u_reg.rf[1][13] ), .QN(_07550_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06530_ ), .Q(\u_reg.rf[1][12] ), .QN(_07551_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06530_ ), .Q(\u_reg.rf[1][29] ), .QN(_07552_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06530_ ), .Q(\u_reg.rf[1][11] ), .QN(_07553_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06530_ ), .Q(\u_reg.rf[1][10] ), .QN(_07554_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06530_ ), .Q(\u_reg.rf[1][9] ), .QN(_07555_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06530_ ), .Q(\u_reg.rf[1][8] ), .QN(_07556_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06530_ ), .Q(\u_reg.rf[1][7] ), .QN(_07557_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06530_ ), .Q(\u_reg.rf[1][6] ), .QN(_07558_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06530_ ), .Q(\u_reg.rf[1][5] ), .QN(_07559_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06530_ ), .Q(\u_reg.rf[1][4] ), .QN(_07560_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06530_ ), .Q(\u_reg.rf[1][3] ), .QN(_07561_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06530_ ), .Q(\u_reg.rf[1][2] ), .QN(_07562_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06530_ ), .Q(\u_reg.rf[1][28] ), .QN(_07563_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06530_ ), .Q(\u_reg.rf[1][1] ), .QN(_07564_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06530_ ), .Q(\u_reg.rf[1][0] ), .QN(_07565_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06530_ ), .Q(\u_reg.rf[1][27] ), .QN(_07566_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06530_ ), .Q(\u_reg.rf[1][26] ), .QN(_07567_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06530_ ), .Q(\u_reg.rf[1][25] ), .QN(_07568_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06530_ ), .Q(\u_reg.rf[1][24] ), .QN(_07569_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06530_ ), .Q(\u_reg.rf[1][23] ), .QN(_07570_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06530_ ), .Q(\u_reg.rf[1][22] ), .QN(_07571_ ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06529_ ), .Q(\u_reg.rf[2][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06529_ ), .Q(\u_reg.rf[2][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06529_ ), .Q(\u_reg.rf[2][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06529_ ), .Q(\u_reg.rf[2][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06529_ ), .Q(\u_reg.rf[2][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06529_ ), .Q(\u_reg.rf[2][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06529_ ), .Q(\u_reg.rf[2][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06529_ ), .Q(\u_reg.rf[2][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06529_ ), .Q(\u_reg.rf[2][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06529_ ), .Q(\u_reg.rf[2][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06529_ ), .Q(\u_reg.rf[2][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06529_ ), .Q(\u_reg.rf[2][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06529_ ), .Q(\u_reg.rf[2][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06529_ ), .Q(\u_reg.rf[2][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06529_ ), .Q(\u_reg.rf[2][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06529_ ), .Q(\u_reg.rf[2][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06529_ ), .Q(\u_reg.rf[2][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06529_ ), .Q(\u_reg.rf[2][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06529_ ), .Q(\u_reg.rf[2][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06529_ ), .Q(\u_reg.rf[2][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06529_ ), .Q(\u_reg.rf[2][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06529_ ), .Q(\u_reg.rf[2][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06529_ ), .Q(\u_reg.rf[2][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06529_ ), .Q(\u_reg.rf[2][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06529_ ), .Q(\u_reg.rf[2][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06529_ ), .Q(\u_reg.rf[2][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06529_ ), .Q(\u_reg.rf[2][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06529_ ), .Q(\u_reg.rf[2][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06529_ ), .Q(\u_reg.rf[2][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06529_ ), .Q(\u_reg.rf[2][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06529_ ), .Q(\u_reg.rf[2][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06529_ ), .Q(\u_reg.rf[2][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06528_ ), .Q(\u_reg.rf[3][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06528_ ), .Q(\u_reg.rf[3][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06528_ ), .Q(\u_reg.rf[3][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06528_ ), .Q(\u_reg.rf[3][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06528_ ), .Q(\u_reg.rf[3][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06528_ ), .Q(\u_reg.rf[3][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06528_ ), .Q(\u_reg.rf[3][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06528_ ), .Q(\u_reg.rf[3][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06528_ ), .Q(\u_reg.rf[3][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06528_ ), .Q(\u_reg.rf[3][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06528_ ), .Q(\u_reg.rf[3][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06528_ ), .Q(\u_reg.rf[3][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06528_ ), .Q(\u_reg.rf[3][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06528_ ), .Q(\u_reg.rf[3][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06528_ ), .Q(\u_reg.rf[3][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06528_ ), .Q(\u_reg.rf[3][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06528_ ), .Q(\u_reg.rf[3][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06528_ ), .Q(\u_reg.rf[3][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06528_ ), .Q(\u_reg.rf[3][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06528_ ), .Q(\u_reg.rf[3][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06528_ ), .Q(\u_reg.rf[3][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06528_ ), .Q(\u_reg.rf[3][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06528_ ), .Q(\u_reg.rf[3][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06528_ ), .Q(\u_reg.rf[3][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06528_ ), .Q(\u_reg.rf[3][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06528_ ), .Q(\u_reg.rf[3][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06528_ ), .Q(\u_reg.rf[3][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06528_ ), .Q(\u_reg.rf[3][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06528_ ), .Q(\u_reg.rf[3][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06528_ ), .Q(\u_reg.rf[3][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06528_ ), .Q(\u_reg.rf[3][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06528_ ), .Q(\u_reg.rf[3][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06527_ ), .Q(\u_reg.rf[4][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06527_ ), .Q(\u_reg.rf[4][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06527_ ), .Q(\u_reg.rf[4][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06527_ ), .Q(\u_reg.rf[4][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06527_ ), .Q(\u_reg.rf[4][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06527_ ), .Q(\u_reg.rf[4][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06527_ ), .Q(\u_reg.rf[4][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06527_ ), .Q(\u_reg.rf[4][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06527_ ), .Q(\u_reg.rf[4][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06527_ ), .Q(\u_reg.rf[4][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06527_ ), .Q(\u_reg.rf[4][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06527_ ), .Q(\u_reg.rf[4][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06527_ ), .Q(\u_reg.rf[4][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06527_ ), .Q(\u_reg.rf[4][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06527_ ), .Q(\u_reg.rf[4][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06527_ ), .Q(\u_reg.rf[4][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06527_ ), .Q(\u_reg.rf[4][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06527_ ), .Q(\u_reg.rf[4][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06527_ ), .Q(\u_reg.rf[4][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06527_ ), .Q(\u_reg.rf[4][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06527_ ), .Q(\u_reg.rf[4][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06527_ ), .Q(\u_reg.rf[4][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06527_ ), .Q(\u_reg.rf[4][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06527_ ), .Q(\u_reg.rf[4][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06527_ ), .Q(\u_reg.rf[4][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06527_ ), .Q(\u_reg.rf[4][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06527_ ), .Q(\u_reg.rf[4][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06527_ ), .Q(\u_reg.rf[4][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06527_ ), .Q(\u_reg.rf[4][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06527_ ), .Q(\u_reg.rf[4][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06527_ ), .Q(\u_reg.rf[4][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06527_ ), .Q(\u_reg.rf[4][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06526_ ), .Q(\u_reg.rf[5][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06526_ ), .Q(\u_reg.rf[5][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06526_ ), .Q(\u_reg.rf[5][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06526_ ), .Q(\u_reg.rf[5][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06526_ ), .Q(\u_reg.rf[5][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06526_ ), .Q(\u_reg.rf[5][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06526_ ), .Q(\u_reg.rf[5][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06526_ ), .Q(\u_reg.rf[5][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06526_ ), .Q(\u_reg.rf[5][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06526_ ), .Q(\u_reg.rf[5][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06526_ ), .Q(\u_reg.rf[5][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06526_ ), .Q(\u_reg.rf[5][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06526_ ), .Q(\u_reg.rf[5][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06526_ ), .Q(\u_reg.rf[5][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06526_ ), .Q(\u_reg.rf[5][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06526_ ), .Q(\u_reg.rf[5][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06526_ ), .Q(\u_reg.rf[5][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06526_ ), .Q(\u_reg.rf[5][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06526_ ), .Q(\u_reg.rf[5][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06526_ ), .Q(\u_reg.rf[5][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06526_ ), .Q(\u_reg.rf[5][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06526_ ), .Q(\u_reg.rf[5][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06526_ ), .Q(\u_reg.rf[5][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06526_ ), .Q(\u_reg.rf[5][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06526_ ), .Q(\u_reg.rf[5][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06526_ ), .Q(\u_reg.rf[5][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06526_ ), .Q(\u_reg.rf[5][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06526_ ), .Q(\u_reg.rf[5][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06526_ ), .Q(\u_reg.rf[5][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06526_ ), .Q(\u_reg.rf[5][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06526_ ), .Q(\u_reg.rf[5][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06526_ ), .Q(\u_reg.rf[5][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06525_ ), .Q(\u_reg.rf[6][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06525_ ), .Q(\u_reg.rf[6][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06525_ ), .Q(\u_reg.rf[6][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06525_ ), .Q(\u_reg.rf[6][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06525_ ), .Q(\u_reg.rf[6][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06525_ ), .Q(\u_reg.rf[6][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06525_ ), .Q(\u_reg.rf[6][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06525_ ), .Q(\u_reg.rf[6][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06525_ ), .Q(\u_reg.rf[6][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06525_ ), .Q(\u_reg.rf[6][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06525_ ), .Q(\u_reg.rf[6][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06525_ ), .Q(\u_reg.rf[6][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06525_ ), .Q(\u_reg.rf[6][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06525_ ), .Q(\u_reg.rf[6][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06525_ ), .Q(\u_reg.rf[6][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06525_ ), .Q(\u_reg.rf[6][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06525_ ), .Q(\u_reg.rf[6][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06525_ ), .Q(\u_reg.rf[6][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06525_ ), .Q(\u_reg.rf[6][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06525_ ), .Q(\u_reg.rf[6][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06525_ ), .Q(\u_reg.rf[6][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06525_ ), .Q(\u_reg.rf[6][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06525_ ), .Q(\u_reg.rf[6][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06525_ ), .Q(\u_reg.rf[6][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06525_ ), .Q(\u_reg.rf[6][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06525_ ), .Q(\u_reg.rf[6][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06525_ ), .Q(\u_reg.rf[6][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06525_ ), .Q(\u_reg.rf[6][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06525_ ), .Q(\u_reg.rf[6][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06525_ ), .Q(\u_reg.rf[6][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06525_ ), .Q(\u_reg.rf[6][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06525_ ), .Q(\u_reg.rf[6][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06524_ ), .Q(\u_reg.rf[7][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06524_ ), .Q(\u_reg.rf[7][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06524_ ), .Q(\u_reg.rf[7][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06524_ ), .Q(\u_reg.rf[7][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06524_ ), .Q(\u_reg.rf[7][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06524_ ), .Q(\u_reg.rf[7][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06524_ ), .Q(\u_reg.rf[7][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06524_ ), .Q(\u_reg.rf[7][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06524_ ), .Q(\u_reg.rf[7][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06524_ ), .Q(\u_reg.rf[7][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06524_ ), .Q(\u_reg.rf[7][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06524_ ), .Q(\u_reg.rf[7][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06524_ ), .Q(\u_reg.rf[7][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06524_ ), .Q(\u_reg.rf[7][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06524_ ), .Q(\u_reg.rf[7][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06524_ ), .Q(\u_reg.rf[7][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06524_ ), .Q(\u_reg.rf[7][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06524_ ), .Q(\u_reg.rf[7][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06524_ ), .Q(\u_reg.rf[7][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06524_ ), .Q(\u_reg.rf[7][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06524_ ), .Q(\u_reg.rf[7][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06524_ ), .Q(\u_reg.rf[7][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06524_ ), .Q(\u_reg.rf[7][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06524_ ), .Q(\u_reg.rf[7][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06524_ ), .Q(\u_reg.rf[7][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06524_ ), .Q(\u_reg.rf[7][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06524_ ), .Q(\u_reg.rf[7][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06524_ ), .Q(\u_reg.rf[7][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06524_ ), .Q(\u_reg.rf[7][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06524_ ), .Q(\u_reg.rf[7][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06524_ ), .Q(\u_reg.rf[7][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06524_ ), .Q(\u_reg.rf[7][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06523_ ), .Q(\u_reg.rf[8][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06523_ ), .Q(\u_reg.rf[8][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06523_ ), .Q(\u_reg.rf[8][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06523_ ), .Q(\u_reg.rf[8][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06523_ ), .Q(\u_reg.rf[8][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06523_ ), .Q(\u_reg.rf[8][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06523_ ), .Q(\u_reg.rf[8][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06523_ ), .Q(\u_reg.rf[8][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06523_ ), .Q(\u_reg.rf[8][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06523_ ), .Q(\u_reg.rf[8][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06523_ ), .Q(\u_reg.rf[8][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06523_ ), .Q(\u_reg.rf[8][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06523_ ), .Q(\u_reg.rf[8][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06523_ ), .Q(\u_reg.rf[8][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06523_ ), .Q(\u_reg.rf[8][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06523_ ), .Q(\u_reg.rf[8][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06523_ ), .Q(\u_reg.rf[8][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06523_ ), .Q(\u_reg.rf[8][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06523_ ), .Q(\u_reg.rf[8][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06523_ ), .Q(\u_reg.rf[8][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06523_ ), .Q(\u_reg.rf[8][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06523_ ), .Q(\u_reg.rf[8][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06523_ ), .Q(\u_reg.rf[8][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06523_ ), .Q(\u_reg.rf[8][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06523_ ), .Q(\u_reg.rf[8][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06523_ ), .Q(\u_reg.rf[8][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06523_ ), .Q(\u_reg.rf[8][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06523_ ), .Q(\u_reg.rf[8][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06523_ ), .Q(\u_reg.rf[8][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06523_ ), .Q(\u_reg.rf[8][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06523_ ), .Q(\u_reg.rf[8][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06523_ ), .Q(\u_reg.rf[8][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q ( .D(\ar_data[31] ), .CK(_06522_ ), .Q(\u_reg.rf[9][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_1 ( .D(\ar_data[30] ), .CK(_06522_ ), .Q(\u_reg.rf[9][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_10 ( .D(\ar_data[21] ), .CK(_06522_ ), .Q(\u_reg.rf[9][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_11 ( .D(\ar_data[20] ), .CK(_06522_ ), .Q(\u_reg.rf[9][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_12 ( .D(\ar_data[19] ), .CK(_06522_ ), .Q(\u_reg.rf[9][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_13 ( .D(\ar_data[18] ), .CK(_06522_ ), .Q(\u_reg.rf[9][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_14 ( .D(\ar_data[17] ), .CK(_06522_ ), .Q(\u_reg.rf[9][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_15 ( .D(\ar_data[16] ), .CK(_06522_ ), .Q(\u_reg.rf[9][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_16 ( .D(\ar_data[15] ), .CK(_06522_ ), .Q(\u_reg.rf[9][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_17 ( .D(\ar_data[14] ), .CK(_06522_ ), .Q(\u_reg.rf[9][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_18 ( .D(\ar_data[13] ), .CK(_06522_ ), .Q(\u_reg.rf[9][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_19 ( .D(\ar_data[12] ), .CK(_06522_ ), .Q(\u_reg.rf[9][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_2 ( .D(\ar_data[29] ), .CK(_06522_ ), .Q(\u_reg.rf[9][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_20 ( .D(\ar_data[11] ), .CK(_06522_ ), .Q(\u_reg.rf[9][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_21 ( .D(\ar_data[10] ), .CK(_06522_ ), .Q(\u_reg.rf[9][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_22 ( .D(\ar_data[9] ), .CK(_06522_ ), .Q(\u_reg.rf[9][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_23 ( .D(\ar_data[8] ), .CK(_06522_ ), .Q(\u_reg.rf[9][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_24 ( .D(\ar_data[7] ), .CK(_06522_ ), .Q(\u_reg.rf[9][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_25 ( .D(\ar_data[6] ), .CK(_06522_ ), .Q(\u_reg.rf[9][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_26 ( .D(\ar_data[5] ), .CK(_06522_ ), .Q(\u_reg.rf[9][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_27 ( .D(\ar_data[4] ), .CK(_06522_ ), .Q(\u_reg.rf[9][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_28 ( .D(\ar_data[3] ), .CK(_06522_ ), .Q(\u_reg.rf[9][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_29 ( .D(\ar_data[2] ), .CK(_06522_ ), .Q(\u_reg.rf[9][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_3 ( .D(\ar_data[28] ), .CK(_06522_ ), .Q(\u_reg.rf[9][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_30 ( .D(\ar_data[1] ), .CK(_06522_ ), .Q(\u_reg.rf[9][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_31 ( .D(\ar_data[0] ), .CK(_06522_ ), .Q(\u_reg.rf[9][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_4 ( .D(\ar_data[27] ), .CK(_06522_ ), .Q(\u_reg.rf[9][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_5 ( .D(\ar_data[26] ), .CK(_06522_ ), .Q(\u_reg.rf[9][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_6 ( .D(\ar_data[25] ), .CK(_06522_ ), .Q(\u_reg.rf[9][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_7 ( .D(\ar_data[24] ), .CK(_06522_ ), .Q(\u_reg.rf[9][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_8 ( .D(\ar_data[23] ), .CK(_06522_ ), .Q(\u_reg.rf[9][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_9 ( .D(\ar_data[22] ), .CK(_06522_ ), .Q(\u_reg.rf[9][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(ea_err ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\fc_addr[2] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\fc_addr[2] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\fc_addr[3] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\fc_addr[3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\fc_addr[4] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\u_arbiter.rvalid ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\u_arbiter.rvalid ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\u_exu.alu_p2[0] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\u_exu.alu_p2[0] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\u_exu.alu_p2[1] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\u_exu.alu_p2[1] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\u_exu.alu_p2[2] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\u_exu.alu_p2[2] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\u_exu.alu_p2[3] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\u_idu.imm_auipc_lui[15] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\u_idu.imm_auipc_lui[20] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\u_idu.imm_auipc_lui[21] ), .Z(fanout_net_23 ) );

endmodule
