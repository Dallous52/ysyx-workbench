// `include "tpdef.vh" 

// module top(
//     input [31:0] inst,
//     output [31:0] pc
// );

//     reg [31:0] rgst [31:0];
    
    

// endmodule

module top(
    input a,
    input b,
    output f
);
    assign f = a ^ b;
endmodule
