//Generate the verilog at 2025-10-20T10:28:17 by iSTA.
module ysyx_25040111 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire de_ard_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire ea_err ;
wire ea_rsign ;
wire exe_valid ;
wire exu_valid ;
wire flush_$_OR__Y_B ;
wire icah_ready ;
wire icah_valid ;
wire idu_ready ;
wire ifu_ready ;
wire io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_B ;
wire io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_B ;
wire io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_B ;
wire io_master_araddr_$_NOT__Y_5_A_$_MUX__Y_A ;
wire io_master_araddr_$_NOT__Y_5_A_$_MUX__Y_B ;
wire io_master_bvalid_$_OR__B_Y ;
wire \u_arbiter.rsign ;
wire \u_arbiter.rvalid ;
wire \u_arbiter.rvalid_$_SDFFE_PP0P__Q_E ;
wire \u_arbiter.working ;
wire \u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ;
wire \u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_AND__A_Y ;
wire \u_arbiter.working_$_SDFFE_PP0P__Q_E ;
wire \u_arbiter.wvalid ;
wire \u_arbiter.wvalid_$_SDFFE_PP0P__Q_E ;
wire \u_csr.csr[0][0] ;
wire \u_csr.csr[0][10] ;
wire \u_csr.csr[0][11] ;
wire \u_csr.csr[0][12] ;
wire \u_csr.csr[0][13] ;
wire \u_csr.csr[0][14] ;
wire \u_csr.csr[0][15] ;
wire \u_csr.csr[0][16] ;
wire \u_csr.csr[0][17] ;
wire \u_csr.csr[0][18] ;
wire \u_csr.csr[0][19] ;
wire \u_csr.csr[0][1] ;
wire \u_csr.csr[0][20] ;
wire \u_csr.csr[0][21] ;
wire \u_csr.csr[0][22] ;
wire \u_csr.csr[0][23] ;
wire \u_csr.csr[0][24] ;
wire \u_csr.csr[0][25] ;
wire \u_csr.csr[0][26] ;
wire \u_csr.csr[0][27] ;
wire \u_csr.csr[0][28] ;
wire \u_csr.csr[0][29] ;
wire \u_csr.csr[0][2] ;
wire \u_csr.csr[0][30] ;
wire \u_csr.csr[0][31] ;
wire \u_csr.csr[0][3] ;
wire \u_csr.csr[0][4] ;
wire \u_csr.csr[0][5] ;
wire \u_csr.csr[0][6] ;
wire \u_csr.csr[0][7] ;
wire \u_csr.csr[0][8] ;
wire \u_csr.csr[0][9] ;
wire \u_csr.csr[1][0] ;
wire \u_csr.csr[1][10] ;
wire \u_csr.csr[1][11] ;
wire \u_csr.csr[1][12] ;
wire \u_csr.csr[1][13] ;
wire \u_csr.csr[1][14] ;
wire \u_csr.csr[1][15] ;
wire \u_csr.csr[1][16] ;
wire \u_csr.csr[1][17] ;
wire \u_csr.csr[1][18] ;
wire \u_csr.csr[1][19] ;
wire \u_csr.csr[1][1] ;
wire \u_csr.csr[1][20] ;
wire \u_csr.csr[1][21] ;
wire \u_csr.csr[1][22] ;
wire \u_csr.csr[1][23] ;
wire \u_csr.csr[1][24] ;
wire \u_csr.csr[1][25] ;
wire \u_csr.csr[1][26] ;
wire \u_csr.csr[1][27] ;
wire \u_csr.csr[1][28] ;
wire \u_csr.csr[1][29] ;
wire \u_csr.csr[1][2] ;
wire \u_csr.csr[1][30] ;
wire \u_csr.csr[1][31] ;
wire \u_csr.csr[1][3] ;
wire \u_csr.csr[1][4] ;
wire \u_csr.csr[1][5] ;
wire \u_csr.csr[1][6] ;
wire \u_csr.csr[1][7] ;
wire \u_csr.csr[1][8] ;
wire \u_csr.csr[1][9] ;
wire \u_csr.csr[2][0] ;
wire \u_csr.csr[2][10] ;
wire \u_csr.csr[2][11] ;
wire \u_csr.csr[2][12] ;
wire \u_csr.csr[2][13] ;
wire \u_csr.csr[2][14] ;
wire \u_csr.csr[2][15] ;
wire \u_csr.csr[2][16] ;
wire \u_csr.csr[2][17] ;
wire \u_csr.csr[2][18] ;
wire \u_csr.csr[2][19] ;
wire \u_csr.csr[2][1] ;
wire \u_csr.csr[2][20] ;
wire \u_csr.csr[2][21] ;
wire \u_csr.csr[2][22] ;
wire \u_csr.csr[2][23] ;
wire \u_csr.csr[2][24] ;
wire \u_csr.csr[2][25] ;
wire \u_csr.csr[2][26] ;
wire \u_csr.csr[2][27] ;
wire \u_csr.csr[2][28] ;
wire \u_csr.csr[2][29] ;
wire \u_csr.csr[2][2] ;
wire \u_csr.csr[2][30] ;
wire \u_csr.csr[2][31] ;
wire \u_csr.csr[2][3] ;
wire \u_csr.csr[2][4] ;
wire \u_csr.csr[2][5] ;
wire \u_csr.csr[2][6] ;
wire \u_csr.csr[2][7] ;
wire \u_csr.csr[2][8] ;
wire \u_csr.csr[2][9] ;
wire \u_csr.csr[3][0] ;
wire \u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y ;
wire \u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire \u_exu.alu_p2_$_SDFFE_PP0P__Q_E ;
wire \u_exu.exe_end_$_ANDNOT__B_Y ;
wire \u_exu.exe_end_$_SDFFE_PP0P__Q_E ;
wire \u_exu.exe_start ;
wire \u_exu.exe_start_$_SDFFE_PP0P__Q_E ;
wire \u_exu.jmpc_ok ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_1_B ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_B ;
wire \u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ;
wire \u_exu.opt_$_NOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B ;
wire \u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ;
wire \u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ;
wire \u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B_$_MUX__B_A_$_NAND__Y_B ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ;
wire \u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_Y_$_MUX__B_A_$_NOR__Y_A_$_ANDNOT__Y_B ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_1_Y_$_AND__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \u_icache.caddr_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ;
wire \u_icache.caddr_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_MUX__B_A ;
wire \u_icache.caddr_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ;
wire \u_icache.caddr_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_MUX__B_A ;
wire \u_icache.caddr_$_SDFFE_PP0P__Q_29_D_$_MUX__B_A ;
wire \u_icache.caddr_$_SDFFE_PP0P__Q_E ;
wire \u_icache.cblocks[0][0] ;
wire \u_icache.cblocks[0][10] ;
wire \u_icache.cblocks[0][11] ;
wire \u_icache.cblocks[0][12] ;
wire \u_icache.cblocks[0][13] ;
wire \u_icache.cblocks[0][14] ;
wire \u_icache.cblocks[0][15] ;
wire \u_icache.cblocks[0][16] ;
wire \u_icache.cblocks[0][17] ;
wire \u_icache.cblocks[0][18] ;
wire \u_icache.cblocks[0][19] ;
wire \u_icache.cblocks[0][1] ;
wire \u_icache.cblocks[0][20] ;
wire \u_icache.cblocks[0][21] ;
wire \u_icache.cblocks[0][22] ;
wire \u_icache.cblocks[0][23] ;
wire \u_icache.cblocks[0][24] ;
wire \u_icache.cblocks[0][25] ;
wire \u_icache.cblocks[0][26] ;
wire \u_icache.cblocks[0][27] ;
wire \u_icache.cblocks[0][28] ;
wire \u_icache.cblocks[0][29] ;
wire \u_icache.cblocks[0][2] ;
wire \u_icache.cblocks[0][30] ;
wire \u_icache.cblocks[0][31] ;
wire \u_icache.cblocks[0][3] ;
wire \u_icache.cblocks[0][4] ;
wire \u_icache.cblocks[0][5] ;
wire \u_icache.cblocks[0][6] ;
wire \u_icache.cblocks[0][7] ;
wire \u_icache.cblocks[0][8] ;
wire \u_icache.cblocks[0][9] ;
wire \u_icache.cblocks[1][0] ;
wire \u_icache.cblocks[1][10] ;
wire \u_icache.cblocks[1][11] ;
wire \u_icache.cblocks[1][12] ;
wire \u_icache.cblocks[1][13] ;
wire \u_icache.cblocks[1][14] ;
wire \u_icache.cblocks[1][15] ;
wire \u_icache.cblocks[1][16] ;
wire \u_icache.cblocks[1][17] ;
wire \u_icache.cblocks[1][18] ;
wire \u_icache.cblocks[1][19] ;
wire \u_icache.cblocks[1][1] ;
wire \u_icache.cblocks[1][20] ;
wire \u_icache.cblocks[1][21] ;
wire \u_icache.cblocks[1][22] ;
wire \u_icache.cblocks[1][23] ;
wire \u_icache.cblocks[1][24] ;
wire \u_icache.cblocks[1][25] ;
wire \u_icache.cblocks[1][26] ;
wire \u_icache.cblocks[1][27] ;
wire \u_icache.cblocks[1][28] ;
wire \u_icache.cblocks[1][29] ;
wire \u_icache.cblocks[1][2] ;
wire \u_icache.cblocks[1][30] ;
wire \u_icache.cblocks[1][31] ;
wire \u_icache.cblocks[1][3] ;
wire \u_icache.cblocks[1][4] ;
wire \u_icache.cblocks[1][5] ;
wire \u_icache.cblocks[1][6] ;
wire \u_icache.cblocks[1][7] ;
wire \u_icache.cblocks[1][8] ;
wire \u_icache.cblocks[1][9] ;
wire \u_icache.cblocks[2][0] ;
wire \u_icache.cblocks[2][10] ;
wire \u_icache.cblocks[2][11] ;
wire \u_icache.cblocks[2][12] ;
wire \u_icache.cblocks[2][13] ;
wire \u_icache.cblocks[2][14] ;
wire \u_icache.cblocks[2][15] ;
wire \u_icache.cblocks[2][16] ;
wire \u_icache.cblocks[2][17] ;
wire \u_icache.cblocks[2][18] ;
wire \u_icache.cblocks[2][19] ;
wire \u_icache.cblocks[2][1] ;
wire \u_icache.cblocks[2][20] ;
wire \u_icache.cblocks[2][21] ;
wire \u_icache.cblocks[2][22] ;
wire \u_icache.cblocks[2][23] ;
wire \u_icache.cblocks[2][24] ;
wire \u_icache.cblocks[2][25] ;
wire \u_icache.cblocks[2][26] ;
wire \u_icache.cblocks[2][27] ;
wire \u_icache.cblocks[2][28] ;
wire \u_icache.cblocks[2][29] ;
wire \u_icache.cblocks[2][2] ;
wire \u_icache.cblocks[2][30] ;
wire \u_icache.cblocks[2][31] ;
wire \u_icache.cblocks[2][3] ;
wire \u_icache.cblocks[2][4] ;
wire \u_icache.cblocks[2][5] ;
wire \u_icache.cblocks[2][6] ;
wire \u_icache.cblocks[2][7] ;
wire \u_icache.cblocks[2][8] ;
wire \u_icache.cblocks[2][9] ;
wire \u_icache.cblocks[3][0] ;
wire \u_icache.cblocks[3][10] ;
wire \u_icache.cblocks[3][11] ;
wire \u_icache.cblocks[3][12] ;
wire \u_icache.cblocks[3][13] ;
wire \u_icache.cblocks[3][14] ;
wire \u_icache.cblocks[3][15] ;
wire \u_icache.cblocks[3][16] ;
wire \u_icache.cblocks[3][17] ;
wire \u_icache.cblocks[3][18] ;
wire \u_icache.cblocks[3][19] ;
wire \u_icache.cblocks[3][1] ;
wire \u_icache.cblocks[3][20] ;
wire \u_icache.cblocks[3][21] ;
wire \u_icache.cblocks[3][22] ;
wire \u_icache.cblocks[3][23] ;
wire \u_icache.cblocks[3][24] ;
wire \u_icache.cblocks[3][25] ;
wire \u_icache.cblocks[3][26] ;
wire \u_icache.cblocks[3][27] ;
wire \u_icache.cblocks[3][28] ;
wire \u_icache.cblocks[3][29] ;
wire \u_icache.cblocks[3][2] ;
wire \u_icache.cblocks[3][30] ;
wire \u_icache.cblocks[3][31] ;
wire \u_icache.cblocks[3][3] ;
wire \u_icache.cblocks[3][4] ;
wire \u_icache.cblocks[3][5] ;
wire \u_icache.cblocks[3][6] ;
wire \u_icache.cblocks[3][7] ;
wire \u_icache.cblocks[3][8] ;
wire \u_icache.cblocks[3][9] ;
wire \u_icache.cblocks[4][0] ;
wire \u_icache.cblocks[4][10] ;
wire \u_icache.cblocks[4][11] ;
wire \u_icache.cblocks[4][12] ;
wire \u_icache.cblocks[4][13] ;
wire \u_icache.cblocks[4][14] ;
wire \u_icache.cblocks[4][15] ;
wire \u_icache.cblocks[4][16] ;
wire \u_icache.cblocks[4][17] ;
wire \u_icache.cblocks[4][18] ;
wire \u_icache.cblocks[4][19] ;
wire \u_icache.cblocks[4][1] ;
wire \u_icache.cblocks[4][20] ;
wire \u_icache.cblocks[4][21] ;
wire \u_icache.cblocks[4][22] ;
wire \u_icache.cblocks[4][23] ;
wire \u_icache.cblocks[4][24] ;
wire \u_icache.cblocks[4][25] ;
wire \u_icache.cblocks[4][26] ;
wire \u_icache.cblocks[4][27] ;
wire \u_icache.cblocks[4][28] ;
wire \u_icache.cblocks[4][29] ;
wire \u_icache.cblocks[4][2] ;
wire \u_icache.cblocks[4][30] ;
wire \u_icache.cblocks[4][31] ;
wire \u_icache.cblocks[4][3] ;
wire \u_icache.cblocks[4][4] ;
wire \u_icache.cblocks[4][5] ;
wire \u_icache.cblocks[4][6] ;
wire \u_icache.cblocks[4][7] ;
wire \u_icache.cblocks[4][8] ;
wire \u_icache.cblocks[4][9] ;
wire \u_icache.cblocks[5][0] ;
wire \u_icache.cblocks[5][10] ;
wire \u_icache.cblocks[5][11] ;
wire \u_icache.cblocks[5][12] ;
wire \u_icache.cblocks[5][13] ;
wire \u_icache.cblocks[5][14] ;
wire \u_icache.cblocks[5][15] ;
wire \u_icache.cblocks[5][16] ;
wire \u_icache.cblocks[5][17] ;
wire \u_icache.cblocks[5][18] ;
wire \u_icache.cblocks[5][19] ;
wire \u_icache.cblocks[5][1] ;
wire \u_icache.cblocks[5][20] ;
wire \u_icache.cblocks[5][21] ;
wire \u_icache.cblocks[5][22] ;
wire \u_icache.cblocks[5][23] ;
wire \u_icache.cblocks[5][24] ;
wire \u_icache.cblocks[5][25] ;
wire \u_icache.cblocks[5][26] ;
wire \u_icache.cblocks[5][27] ;
wire \u_icache.cblocks[5][28] ;
wire \u_icache.cblocks[5][29] ;
wire \u_icache.cblocks[5][2] ;
wire \u_icache.cblocks[5][30] ;
wire \u_icache.cblocks[5][31] ;
wire \u_icache.cblocks[5][3] ;
wire \u_icache.cblocks[5][4] ;
wire \u_icache.cblocks[5][5] ;
wire \u_icache.cblocks[5][6] ;
wire \u_icache.cblocks[5][7] ;
wire \u_icache.cblocks[5][8] ;
wire \u_icache.cblocks[5][9] ;
wire \u_icache.cblocks[6][0] ;
wire \u_icache.cblocks[6][10] ;
wire \u_icache.cblocks[6][11] ;
wire \u_icache.cblocks[6][12] ;
wire \u_icache.cblocks[6][13] ;
wire \u_icache.cblocks[6][14] ;
wire \u_icache.cblocks[6][15] ;
wire \u_icache.cblocks[6][16] ;
wire \u_icache.cblocks[6][17] ;
wire \u_icache.cblocks[6][18] ;
wire \u_icache.cblocks[6][19] ;
wire \u_icache.cblocks[6][1] ;
wire \u_icache.cblocks[6][20] ;
wire \u_icache.cblocks[6][21] ;
wire \u_icache.cblocks[6][22] ;
wire \u_icache.cblocks[6][23] ;
wire \u_icache.cblocks[6][24] ;
wire \u_icache.cblocks[6][25] ;
wire \u_icache.cblocks[6][26] ;
wire \u_icache.cblocks[6][27] ;
wire \u_icache.cblocks[6][28] ;
wire \u_icache.cblocks[6][29] ;
wire \u_icache.cblocks[6][2] ;
wire \u_icache.cblocks[6][30] ;
wire \u_icache.cblocks[6][31] ;
wire \u_icache.cblocks[6][3] ;
wire \u_icache.cblocks[6][4] ;
wire \u_icache.cblocks[6][5] ;
wire \u_icache.cblocks[6][6] ;
wire \u_icache.cblocks[6][7] ;
wire \u_icache.cblocks[6][8] ;
wire \u_icache.cblocks[6][9] ;
wire \u_icache.cblocks[7][0] ;
wire \u_icache.cblocks[7][10] ;
wire \u_icache.cblocks[7][11] ;
wire \u_icache.cblocks[7][12] ;
wire \u_icache.cblocks[7][13] ;
wire \u_icache.cblocks[7][14] ;
wire \u_icache.cblocks[7][15] ;
wire \u_icache.cblocks[7][16] ;
wire \u_icache.cblocks[7][17] ;
wire \u_icache.cblocks[7][18] ;
wire \u_icache.cblocks[7][19] ;
wire \u_icache.cblocks[7][1] ;
wire \u_icache.cblocks[7][20] ;
wire \u_icache.cblocks[7][21] ;
wire \u_icache.cblocks[7][22] ;
wire \u_icache.cblocks[7][23] ;
wire \u_icache.cblocks[7][24] ;
wire \u_icache.cblocks[7][25] ;
wire \u_icache.cblocks[7][26] ;
wire \u_icache.cblocks[7][27] ;
wire \u_icache.cblocks[7][28] ;
wire \u_icache.cblocks[7][29] ;
wire \u_icache.cblocks[7][2] ;
wire \u_icache.cblocks[7][30] ;
wire \u_icache.cblocks[7][31] ;
wire \u_icache.cblocks[7][3] ;
wire \u_icache.cblocks[7][4] ;
wire \u_icache.cblocks[7][5] ;
wire \u_icache.cblocks[7][6] ;
wire \u_icache.cblocks[7][7] ;
wire \u_icache.cblocks[7][8] ;
wire \u_icache.cblocks[7][9] ;
wire \u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ;
wire \u_icache.chvalid_$_SDFFE_PP0P__Q_E ;
wire \u_icache.count_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_NOT__A_Y ;
wire \u_icache.count_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_ORNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_OR__B_1_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_OR__B_2_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_OR__B_3_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \u_icache.count_$_SDFFE_PP0P__Q_E ;
wire \u_icache.cready_$_ANDNOT__A_Y ;
wire \u_icache.cready_$_ANDNOT__B_Y_$_OR__B_Y ;
wire \u_icache.ctags[0][0] ;
wire \u_icache.ctags[0][10] ;
wire \u_icache.ctags[0][11] ;
wire \u_icache.ctags[0][12] ;
wire \u_icache.ctags[0][13] ;
wire \u_icache.ctags[0][14] ;
wire \u_icache.ctags[0][15] ;
wire \u_icache.ctags[0][16] ;
wire \u_icache.ctags[0][17] ;
wire \u_icache.ctags[0][18] ;
wire \u_icache.ctags[0][19] ;
wire \u_icache.ctags[0][1] ;
wire \u_icache.ctags[0][20] ;
wire \u_icache.ctags[0][21] ;
wire \u_icache.ctags[0][22] ;
wire \u_icache.ctags[0][23] ;
wire \u_icache.ctags[0][24] ;
wire \u_icache.ctags[0][25] ;
wire \u_icache.ctags[0][26] ;
wire \u_icache.ctags[0][2] ;
wire \u_icache.ctags[0][3] ;
wire \u_icache.ctags[0][4] ;
wire \u_icache.ctags[0][5] ;
wire \u_icache.ctags[0][6] ;
wire \u_icache.ctags[0][7] ;
wire \u_icache.ctags[0][8] ;
wire \u_icache.ctags[0][9] ;
wire \u_icache.ctags[1][0] ;
wire \u_icache.ctags[1][10] ;
wire \u_icache.ctags[1][11] ;
wire \u_icache.ctags[1][12] ;
wire \u_icache.ctags[1][13] ;
wire \u_icache.ctags[1][14] ;
wire \u_icache.ctags[1][15] ;
wire \u_icache.ctags[1][16] ;
wire \u_icache.ctags[1][17] ;
wire \u_icache.ctags[1][18] ;
wire \u_icache.ctags[1][19] ;
wire \u_icache.ctags[1][1] ;
wire \u_icache.ctags[1][20] ;
wire \u_icache.ctags[1][21] ;
wire \u_icache.ctags[1][22] ;
wire \u_icache.ctags[1][23] ;
wire \u_icache.ctags[1][24] ;
wire \u_icache.ctags[1][25] ;
wire \u_icache.ctags[1][26] ;
wire \u_icache.ctags[1][2] ;
wire \u_icache.ctags[1][3] ;
wire \u_icache.ctags[1][4] ;
wire \u_icache.ctags[1][5] ;
wire \u_icache.ctags[1][6] ;
wire \u_icache.ctags[1][7] ;
wire \u_icache.ctags[1][8] ;
wire \u_icache.ctags[1][9] ;
wire \u_icache.cvalids_$_SDFFE_PP0P__Q_E ;
wire \u_icache.ended ;
wire \u_icache.ended_$_SDFFE_PP0P__Q_E ;
wire \u_idu.decode_ok_$_SDFFE_PP0P__Q_E ;
wire \u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ;
wire \u_ifu.inst_ok_$_ANDNOT__A_Y ;
wire \u_ifu.inst_ok_$_SDFFE_PP0P__Q_E ;
wire \u_ifu.jpc_ok ;
wire \u_ifu.jpc_ok_$_NOT__A_Y ;
wire \u_ifu.jpc_ok_$_SDFFE_PP0P__Q_E ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_B_$_ANDNOT__B_Y ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_Y ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ;
wire \u_ifu.pc_$_SDFFE_PP0N__Q_28_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \u_ifu.pc_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.arvalid ;
wire \u_lsu.arvalid_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.awvalid_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.reading ;
wire \u_lsu.reading_$_NOR__B_A_$_MUX__Y_A ;
wire \u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ;
wire \u_lsu.reading_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.rvalid ;
wire \u_lsu.rvalid_clint ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_10_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_18_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_26_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_28_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_31_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_39_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_8_A_$_ANDNOT__Y_B ;
wire \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ;
wire \u_lsu.wlast_$_SDFFE_PP0P__Q_E ;
wire \u_lsu.writing ;
wire \u_reg.rf[10][0] ;
wire \u_reg.rf[10][10] ;
wire \u_reg.rf[10][11] ;
wire \u_reg.rf[10][12] ;
wire \u_reg.rf[10][13] ;
wire \u_reg.rf[10][14] ;
wire \u_reg.rf[10][15] ;
wire \u_reg.rf[10][16] ;
wire \u_reg.rf[10][17] ;
wire \u_reg.rf[10][18] ;
wire \u_reg.rf[10][19] ;
wire \u_reg.rf[10][1] ;
wire \u_reg.rf[10][20] ;
wire \u_reg.rf[10][21] ;
wire \u_reg.rf[10][22] ;
wire \u_reg.rf[10][23] ;
wire \u_reg.rf[10][24] ;
wire \u_reg.rf[10][25] ;
wire \u_reg.rf[10][26] ;
wire \u_reg.rf[10][27] ;
wire \u_reg.rf[10][28] ;
wire \u_reg.rf[10][29] ;
wire \u_reg.rf[10][2] ;
wire \u_reg.rf[10][30] ;
wire \u_reg.rf[10][31] ;
wire \u_reg.rf[10][3] ;
wire \u_reg.rf[10][4] ;
wire \u_reg.rf[10][5] ;
wire \u_reg.rf[10][6] ;
wire \u_reg.rf[10][7] ;
wire \u_reg.rf[10][8] ;
wire \u_reg.rf[10][9] ;
wire \u_reg.rf[11][0] ;
wire \u_reg.rf[11][10] ;
wire \u_reg.rf[11][11] ;
wire \u_reg.rf[11][12] ;
wire \u_reg.rf[11][13] ;
wire \u_reg.rf[11][14] ;
wire \u_reg.rf[11][15] ;
wire \u_reg.rf[11][16] ;
wire \u_reg.rf[11][17] ;
wire \u_reg.rf[11][18] ;
wire \u_reg.rf[11][19] ;
wire \u_reg.rf[11][1] ;
wire \u_reg.rf[11][20] ;
wire \u_reg.rf[11][21] ;
wire \u_reg.rf[11][22] ;
wire \u_reg.rf[11][23] ;
wire \u_reg.rf[11][24] ;
wire \u_reg.rf[11][25] ;
wire \u_reg.rf[11][26] ;
wire \u_reg.rf[11][27] ;
wire \u_reg.rf[11][28] ;
wire \u_reg.rf[11][29] ;
wire \u_reg.rf[11][2] ;
wire \u_reg.rf[11][30] ;
wire \u_reg.rf[11][31] ;
wire \u_reg.rf[11][3] ;
wire \u_reg.rf[11][4] ;
wire \u_reg.rf[11][5] ;
wire \u_reg.rf[11][6] ;
wire \u_reg.rf[11][7] ;
wire \u_reg.rf[11][8] ;
wire \u_reg.rf[11][9] ;
wire \u_reg.rf[12][0] ;
wire \u_reg.rf[12][10] ;
wire \u_reg.rf[12][11] ;
wire \u_reg.rf[12][12] ;
wire \u_reg.rf[12][13] ;
wire \u_reg.rf[12][14] ;
wire \u_reg.rf[12][15] ;
wire \u_reg.rf[12][16] ;
wire \u_reg.rf[12][17] ;
wire \u_reg.rf[12][18] ;
wire \u_reg.rf[12][19] ;
wire \u_reg.rf[12][1] ;
wire \u_reg.rf[12][20] ;
wire \u_reg.rf[12][21] ;
wire \u_reg.rf[12][22] ;
wire \u_reg.rf[12][23] ;
wire \u_reg.rf[12][24] ;
wire \u_reg.rf[12][25] ;
wire \u_reg.rf[12][26] ;
wire \u_reg.rf[12][27] ;
wire \u_reg.rf[12][28] ;
wire \u_reg.rf[12][29] ;
wire \u_reg.rf[12][2] ;
wire \u_reg.rf[12][30] ;
wire \u_reg.rf[12][31] ;
wire \u_reg.rf[12][3] ;
wire \u_reg.rf[12][4] ;
wire \u_reg.rf[12][5] ;
wire \u_reg.rf[12][6] ;
wire \u_reg.rf[12][7] ;
wire \u_reg.rf[12][8] ;
wire \u_reg.rf[12][9] ;
wire \u_reg.rf[13][0] ;
wire \u_reg.rf[13][10] ;
wire \u_reg.rf[13][11] ;
wire \u_reg.rf[13][12] ;
wire \u_reg.rf[13][13] ;
wire \u_reg.rf[13][14] ;
wire \u_reg.rf[13][15] ;
wire \u_reg.rf[13][16] ;
wire \u_reg.rf[13][17] ;
wire \u_reg.rf[13][18] ;
wire \u_reg.rf[13][19] ;
wire \u_reg.rf[13][1] ;
wire \u_reg.rf[13][20] ;
wire \u_reg.rf[13][21] ;
wire \u_reg.rf[13][22] ;
wire \u_reg.rf[13][23] ;
wire \u_reg.rf[13][24] ;
wire \u_reg.rf[13][25] ;
wire \u_reg.rf[13][26] ;
wire \u_reg.rf[13][27] ;
wire \u_reg.rf[13][28] ;
wire \u_reg.rf[13][29] ;
wire \u_reg.rf[13][2] ;
wire \u_reg.rf[13][30] ;
wire \u_reg.rf[13][31] ;
wire \u_reg.rf[13][3] ;
wire \u_reg.rf[13][4] ;
wire \u_reg.rf[13][5] ;
wire \u_reg.rf[13][6] ;
wire \u_reg.rf[13][7] ;
wire \u_reg.rf[13][8] ;
wire \u_reg.rf[13][9] ;
wire \u_reg.rf[14][0] ;
wire \u_reg.rf[14][10] ;
wire \u_reg.rf[14][11] ;
wire \u_reg.rf[14][12] ;
wire \u_reg.rf[14][13] ;
wire \u_reg.rf[14][14] ;
wire \u_reg.rf[14][15] ;
wire \u_reg.rf[14][16] ;
wire \u_reg.rf[14][17] ;
wire \u_reg.rf[14][18] ;
wire \u_reg.rf[14][19] ;
wire \u_reg.rf[14][1] ;
wire \u_reg.rf[14][20] ;
wire \u_reg.rf[14][21] ;
wire \u_reg.rf[14][22] ;
wire \u_reg.rf[14][23] ;
wire \u_reg.rf[14][24] ;
wire \u_reg.rf[14][25] ;
wire \u_reg.rf[14][26] ;
wire \u_reg.rf[14][27] ;
wire \u_reg.rf[14][28] ;
wire \u_reg.rf[14][29] ;
wire \u_reg.rf[14][2] ;
wire \u_reg.rf[14][30] ;
wire \u_reg.rf[14][31] ;
wire \u_reg.rf[14][3] ;
wire \u_reg.rf[14][4] ;
wire \u_reg.rf[14][5] ;
wire \u_reg.rf[14][6] ;
wire \u_reg.rf[14][7] ;
wire \u_reg.rf[14][8] ;
wire \u_reg.rf[14][9] ;
wire \u_reg.rf[15][0] ;
wire \u_reg.rf[15][10] ;
wire \u_reg.rf[15][11] ;
wire \u_reg.rf[15][12] ;
wire \u_reg.rf[15][13] ;
wire \u_reg.rf[15][14] ;
wire \u_reg.rf[15][15] ;
wire \u_reg.rf[15][16] ;
wire \u_reg.rf[15][17] ;
wire \u_reg.rf[15][18] ;
wire \u_reg.rf[15][19] ;
wire \u_reg.rf[15][1] ;
wire \u_reg.rf[15][20] ;
wire \u_reg.rf[15][21] ;
wire \u_reg.rf[15][22] ;
wire \u_reg.rf[15][23] ;
wire \u_reg.rf[15][24] ;
wire \u_reg.rf[15][25] ;
wire \u_reg.rf[15][26] ;
wire \u_reg.rf[15][27] ;
wire \u_reg.rf[15][28] ;
wire \u_reg.rf[15][29] ;
wire \u_reg.rf[15][2] ;
wire \u_reg.rf[15][30] ;
wire \u_reg.rf[15][31] ;
wire \u_reg.rf[15][3] ;
wire \u_reg.rf[15][4] ;
wire \u_reg.rf[15][5] ;
wire \u_reg.rf[15][6] ;
wire \u_reg.rf[15][7] ;
wire \u_reg.rf[15][8] ;
wire \u_reg.rf[15][9] ;
wire \u_reg.rf[1][0] ;
wire \u_reg.rf[1][10] ;
wire \u_reg.rf[1][11] ;
wire \u_reg.rf[1][12] ;
wire \u_reg.rf[1][13] ;
wire \u_reg.rf[1][14] ;
wire \u_reg.rf[1][15] ;
wire \u_reg.rf[1][16] ;
wire \u_reg.rf[1][17] ;
wire \u_reg.rf[1][18] ;
wire \u_reg.rf[1][19] ;
wire \u_reg.rf[1][1] ;
wire \u_reg.rf[1][20] ;
wire \u_reg.rf[1][21] ;
wire \u_reg.rf[1][22] ;
wire \u_reg.rf[1][23] ;
wire \u_reg.rf[1][24] ;
wire \u_reg.rf[1][25] ;
wire \u_reg.rf[1][26] ;
wire \u_reg.rf[1][27] ;
wire \u_reg.rf[1][28] ;
wire \u_reg.rf[1][29] ;
wire \u_reg.rf[1][2] ;
wire \u_reg.rf[1][30] ;
wire \u_reg.rf[1][31] ;
wire \u_reg.rf[1][3] ;
wire \u_reg.rf[1][4] ;
wire \u_reg.rf[1][5] ;
wire \u_reg.rf[1][6] ;
wire \u_reg.rf[1][7] ;
wire \u_reg.rf[1][8] ;
wire \u_reg.rf[1][9] ;
wire \u_reg.rf[2][0] ;
wire \u_reg.rf[2][10] ;
wire \u_reg.rf[2][11] ;
wire \u_reg.rf[2][12] ;
wire \u_reg.rf[2][13] ;
wire \u_reg.rf[2][14] ;
wire \u_reg.rf[2][15] ;
wire \u_reg.rf[2][16] ;
wire \u_reg.rf[2][17] ;
wire \u_reg.rf[2][18] ;
wire \u_reg.rf[2][19] ;
wire \u_reg.rf[2][1] ;
wire \u_reg.rf[2][20] ;
wire \u_reg.rf[2][21] ;
wire \u_reg.rf[2][22] ;
wire \u_reg.rf[2][23] ;
wire \u_reg.rf[2][24] ;
wire \u_reg.rf[2][25] ;
wire \u_reg.rf[2][26] ;
wire \u_reg.rf[2][27] ;
wire \u_reg.rf[2][28] ;
wire \u_reg.rf[2][29] ;
wire \u_reg.rf[2][2] ;
wire \u_reg.rf[2][30] ;
wire \u_reg.rf[2][31] ;
wire \u_reg.rf[2][3] ;
wire \u_reg.rf[2][4] ;
wire \u_reg.rf[2][5] ;
wire \u_reg.rf[2][6] ;
wire \u_reg.rf[2][7] ;
wire \u_reg.rf[2][8] ;
wire \u_reg.rf[2][9] ;
wire \u_reg.rf[3][0] ;
wire \u_reg.rf[3][10] ;
wire \u_reg.rf[3][11] ;
wire \u_reg.rf[3][12] ;
wire \u_reg.rf[3][13] ;
wire \u_reg.rf[3][14] ;
wire \u_reg.rf[3][15] ;
wire \u_reg.rf[3][16] ;
wire \u_reg.rf[3][17] ;
wire \u_reg.rf[3][18] ;
wire \u_reg.rf[3][19] ;
wire \u_reg.rf[3][1] ;
wire \u_reg.rf[3][20] ;
wire \u_reg.rf[3][21] ;
wire \u_reg.rf[3][22] ;
wire \u_reg.rf[3][23] ;
wire \u_reg.rf[3][24] ;
wire \u_reg.rf[3][25] ;
wire \u_reg.rf[3][26] ;
wire \u_reg.rf[3][27] ;
wire \u_reg.rf[3][28] ;
wire \u_reg.rf[3][29] ;
wire \u_reg.rf[3][2] ;
wire \u_reg.rf[3][30] ;
wire \u_reg.rf[3][31] ;
wire \u_reg.rf[3][3] ;
wire \u_reg.rf[3][4] ;
wire \u_reg.rf[3][5] ;
wire \u_reg.rf[3][6] ;
wire \u_reg.rf[3][7] ;
wire \u_reg.rf[3][8] ;
wire \u_reg.rf[3][9] ;
wire \u_reg.rf[4][0] ;
wire \u_reg.rf[4][10] ;
wire \u_reg.rf[4][11] ;
wire \u_reg.rf[4][12] ;
wire \u_reg.rf[4][13] ;
wire \u_reg.rf[4][14] ;
wire \u_reg.rf[4][15] ;
wire \u_reg.rf[4][16] ;
wire \u_reg.rf[4][17] ;
wire \u_reg.rf[4][18] ;
wire \u_reg.rf[4][19] ;
wire \u_reg.rf[4][1] ;
wire \u_reg.rf[4][20] ;
wire \u_reg.rf[4][21] ;
wire \u_reg.rf[4][22] ;
wire \u_reg.rf[4][23] ;
wire \u_reg.rf[4][24] ;
wire \u_reg.rf[4][25] ;
wire \u_reg.rf[4][26] ;
wire \u_reg.rf[4][27] ;
wire \u_reg.rf[4][28] ;
wire \u_reg.rf[4][29] ;
wire \u_reg.rf[4][2] ;
wire \u_reg.rf[4][30] ;
wire \u_reg.rf[4][31] ;
wire \u_reg.rf[4][3] ;
wire \u_reg.rf[4][4] ;
wire \u_reg.rf[4][5] ;
wire \u_reg.rf[4][6] ;
wire \u_reg.rf[4][7] ;
wire \u_reg.rf[4][8] ;
wire \u_reg.rf[4][9] ;
wire \u_reg.rf[5][0] ;
wire \u_reg.rf[5][10] ;
wire \u_reg.rf[5][11] ;
wire \u_reg.rf[5][12] ;
wire \u_reg.rf[5][13] ;
wire \u_reg.rf[5][14] ;
wire \u_reg.rf[5][15] ;
wire \u_reg.rf[5][16] ;
wire \u_reg.rf[5][17] ;
wire \u_reg.rf[5][18] ;
wire \u_reg.rf[5][19] ;
wire \u_reg.rf[5][1] ;
wire \u_reg.rf[5][20] ;
wire \u_reg.rf[5][21] ;
wire \u_reg.rf[5][22] ;
wire \u_reg.rf[5][23] ;
wire \u_reg.rf[5][24] ;
wire \u_reg.rf[5][25] ;
wire \u_reg.rf[5][26] ;
wire \u_reg.rf[5][27] ;
wire \u_reg.rf[5][28] ;
wire \u_reg.rf[5][29] ;
wire \u_reg.rf[5][2] ;
wire \u_reg.rf[5][30] ;
wire \u_reg.rf[5][31] ;
wire \u_reg.rf[5][3] ;
wire \u_reg.rf[5][4] ;
wire \u_reg.rf[5][5] ;
wire \u_reg.rf[5][6] ;
wire \u_reg.rf[5][7] ;
wire \u_reg.rf[5][8] ;
wire \u_reg.rf[5][9] ;
wire \u_reg.rf[6][0] ;
wire \u_reg.rf[6][10] ;
wire \u_reg.rf[6][11] ;
wire \u_reg.rf[6][12] ;
wire \u_reg.rf[6][13] ;
wire \u_reg.rf[6][14] ;
wire \u_reg.rf[6][15] ;
wire \u_reg.rf[6][16] ;
wire \u_reg.rf[6][17] ;
wire \u_reg.rf[6][18] ;
wire \u_reg.rf[6][19] ;
wire \u_reg.rf[6][1] ;
wire \u_reg.rf[6][20] ;
wire \u_reg.rf[6][21] ;
wire \u_reg.rf[6][22] ;
wire \u_reg.rf[6][23] ;
wire \u_reg.rf[6][24] ;
wire \u_reg.rf[6][25] ;
wire \u_reg.rf[6][26] ;
wire \u_reg.rf[6][27] ;
wire \u_reg.rf[6][28] ;
wire \u_reg.rf[6][29] ;
wire \u_reg.rf[6][2] ;
wire \u_reg.rf[6][30] ;
wire \u_reg.rf[6][31] ;
wire \u_reg.rf[6][3] ;
wire \u_reg.rf[6][4] ;
wire \u_reg.rf[6][5] ;
wire \u_reg.rf[6][6] ;
wire \u_reg.rf[6][7] ;
wire \u_reg.rf[6][8] ;
wire \u_reg.rf[6][9] ;
wire \u_reg.rf[7][0] ;
wire \u_reg.rf[7][10] ;
wire \u_reg.rf[7][11] ;
wire \u_reg.rf[7][12] ;
wire \u_reg.rf[7][13] ;
wire \u_reg.rf[7][14] ;
wire \u_reg.rf[7][15] ;
wire \u_reg.rf[7][16] ;
wire \u_reg.rf[7][17] ;
wire \u_reg.rf[7][18] ;
wire \u_reg.rf[7][19] ;
wire \u_reg.rf[7][1] ;
wire \u_reg.rf[7][20] ;
wire \u_reg.rf[7][21] ;
wire \u_reg.rf[7][22] ;
wire \u_reg.rf[7][23] ;
wire \u_reg.rf[7][24] ;
wire \u_reg.rf[7][25] ;
wire \u_reg.rf[7][26] ;
wire \u_reg.rf[7][27] ;
wire \u_reg.rf[7][28] ;
wire \u_reg.rf[7][29] ;
wire \u_reg.rf[7][2] ;
wire \u_reg.rf[7][30] ;
wire \u_reg.rf[7][31] ;
wire \u_reg.rf[7][3] ;
wire \u_reg.rf[7][4] ;
wire \u_reg.rf[7][5] ;
wire \u_reg.rf[7][6] ;
wire \u_reg.rf[7][7] ;
wire \u_reg.rf[7][8] ;
wire \u_reg.rf[7][9] ;
wire \u_reg.rf[8][0] ;
wire \u_reg.rf[8][10] ;
wire \u_reg.rf[8][11] ;
wire \u_reg.rf[8][12] ;
wire \u_reg.rf[8][13] ;
wire \u_reg.rf[8][14] ;
wire \u_reg.rf[8][15] ;
wire \u_reg.rf[8][16] ;
wire \u_reg.rf[8][17] ;
wire \u_reg.rf[8][18] ;
wire \u_reg.rf[8][19] ;
wire \u_reg.rf[8][1] ;
wire \u_reg.rf[8][20] ;
wire \u_reg.rf[8][21] ;
wire \u_reg.rf[8][22] ;
wire \u_reg.rf[8][23] ;
wire \u_reg.rf[8][24] ;
wire \u_reg.rf[8][25] ;
wire \u_reg.rf[8][26] ;
wire \u_reg.rf[8][27] ;
wire \u_reg.rf[8][28] ;
wire \u_reg.rf[8][29] ;
wire \u_reg.rf[8][2] ;
wire \u_reg.rf[8][30] ;
wire \u_reg.rf[8][31] ;
wire \u_reg.rf[8][3] ;
wire \u_reg.rf[8][4] ;
wire \u_reg.rf[8][5] ;
wire \u_reg.rf[8][6] ;
wire \u_reg.rf[8][7] ;
wire \u_reg.rf[8][8] ;
wire \u_reg.rf[8][9] ;
wire \u_reg.rf[9][0] ;
wire \u_reg.rf[9][10] ;
wire \u_reg.rf[9][11] ;
wire \u_reg.rf[9][12] ;
wire \u_reg.rf[9][13] ;
wire \u_reg.rf[9][14] ;
wire \u_reg.rf[9][15] ;
wire \u_reg.rf[9][16] ;
wire \u_reg.rf[9][17] ;
wire \u_reg.rf[9][18] ;
wire \u_reg.rf[9][19] ;
wire \u_reg.rf[9][1] ;
wire \u_reg.rf[9][20] ;
wire \u_reg.rf[9][21] ;
wire \u_reg.rf[9][22] ;
wire \u_reg.rf[9][23] ;
wire \u_reg.rf[9][24] ;
wire \u_reg.rf[9][25] ;
wire \u_reg.rf[9][26] ;
wire \u_reg.rf[9][27] ;
wire \u_reg.rf[9][28] ;
wire \u_reg.rf[9][29] ;
wire \u_reg.rf[9][2] ;
wire \u_reg.rf[9][30] ;
wire \u_reg.rf[9][31] ;
wire \u_reg.rf[9][3] ;
wire \u_reg.rf[9][4] ;
wire \u_reg.rf[9][5] ;
wire \u_reg.rf[9][6] ;
wire \u_reg.rf[9][7] ;
wire \u_reg.rf[9][8] ;
wire \u_reg.rf[9][9] ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] ac_data ;
wire [31:0] al_wdata ;
wire [1:0] al_wmask ;
wire [31:0] ar_data ;
wire [31:0] ca_addr ;
wire [31:0] cf_inst ;
wire [31:0] de_pc ;
wire [31:0] ea_addr ;
wire [3:0] ea_ard ;
wire [0:0] ea_errtp ;
wire [1:0] ea_mask ;
wire [31:0] ea_pc ;
wire [31:0] ea_wdata ;
wire [31:0] fc_addr ;
wire [31:0] fd_inst ;
wire [31:0] \u_arbiter.raddr ;
wire [1:0] \u_arbiter.rmask ;
wire [3:0] \u_arbiter.wbaddr ;
wire [11:0] \u_exu.acsrd ;
wire [6:0] \u_exu.alu_ctrl ;
wire [31:0] \u_exu.alu_p1 ;
wire [31:0] \u_exu.alu_p2 ;
wire [31:0] \u_exu.ecsr ;
wire [15:0] \u_exu.eopt ;
wire [15:0] \u_exu.rlock ;
wire [0:0] \u_icache.caddr_$_SDFFE_PP0P__Q_28_D ;
wire [2:0] \u_icache.count ;
wire [1:0] \u_icache.cvalids ;
wire [31:0] \u_idu.imm_auipc_lui ;
wire [11:0] \u_idu.imm_branch ;
wire [6:0] \u_idu.inst ;
wire [7:0] \u_lsu.rcount ;
wire [63:0] \u_lsu.u_clint.mtime ;
wire [0:0] \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D ;

assign \io_master_awid [0] = \io_master_arburst [0] ;
assign \io_master_awid [1] = \io_master_arburst [0] ;
assign \io_master_awid [2] = \io_master_arburst [0] ;
assign \io_master_awid [3] = \io_master_arburst [0] ;
assign \io_master_awlen [0] = \io_master_arburst [0] ;
assign \io_master_awlen [1] = \io_master_arburst [0] ;
assign \io_master_awlen [2] = \io_master_arburst [0] ;
assign \io_master_awlen [3] = \io_master_arburst [0] ;
assign \io_master_awlen [4] = \io_master_arburst [0] ;
assign \io_master_awlen [5] = \io_master_arburst [0] ;
assign \io_master_awlen [6] = \io_master_arburst [0] ;
assign \io_master_awlen [7] = \io_master_arburst [0] ;
assign \io_master_awsize [2] = \io_master_arburst [0] ;
assign \io_master_awburst [0] = \io_master_arburst [0] ;
assign \io_master_awburst [1] = \io_master_arburst [0] ;
assign io_master_wvalid = io_master_wlast ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [1] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [0] ;
assign \io_master_arid [3] = \io_master_arburst [0] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [0] ;
assign \io_master_arlen [2] = \io_master_arburst [0] ;
assign \io_master_arlen [3] = \io_master_arburst [0] ;
assign \io_master_arlen [4] = \io_master_arburst [0] ;
assign \io_master_arlen [5] = \io_master_arburst [0] ;
assign \io_master_arlen [6] = \io_master_arburst [0] ;
assign \io_master_arlen [7] = \io_master_arburst [0] ;
assign \io_master_arsize [2] = \io_master_arburst [0] ;
assign \io_master_arburst [1] = \io_master_arburst [0] ;

INV_X1 _07660_ ( .A(\ea_mask [1] ), .ZN(_00629_ ) );
INV_X1 _07661_ ( .A(\ea_mask [0] ), .ZN(_00630_ ) );
AOI21_X1 _07662_ ( .A(\u_exu.eopt [15] ), .B1(_00629_ ), .B2(_00630_ ), .ZN(_00631_ ) );
OR2_X1 _07663_ ( .A1(_00631_ ), .A2(fanout_net_5 ), .ZN(_00632_ ) );
AND2_X1 _07664_ ( .A1(_00632_ ), .A2(icah_valid ), .ZN(_00633_ ) );
INV_X32 _07665_ ( .A(\u_arbiter.working ), .ZN(_00634_ ) );
BUF_X16 _07666_ ( .A(_00634_ ), .Z(_00635_ ) );
NAND2_X1 _07667_ ( .A1(_00635_ ), .A2(exu_valid ), .ZN(_00636_ ) );
NOR2_X1 _07668_ ( .A1(_00633_ ), .A2(_00636_ ), .ZN(_00637_ ) );
AND2_X2 _07669_ ( .A1(_00637_ ), .A2(fanout_net_5 ), .ZN(_00638_ ) );
INV_X2 _07670_ ( .A(_00638_ ), .ZN(_00639_ ) );
BUF_X4 _07671_ ( .A(_00639_ ), .Z(_00640_ ) );
NOR2_X1 _07672_ ( .A1(\u_idu.imm_auipc_lui [28] ), .A2(\u_idu.imm_auipc_lui [29] ), .ZN(_00641_ ) );
NOR2_X1 _07673_ ( .A1(\u_idu.imm_auipc_lui [27] ), .A2(\u_idu.imm_auipc_lui [26] ), .ZN(_00642_ ) );
AND2_X1 _07674_ ( .A1(_00641_ ), .A2(_00642_ ), .ZN(_00643_ ) );
NOR2_X1 _07675_ ( .A1(\u_idu.imm_auipc_lui [31] ), .A2(\u_idu.imm_auipc_lui [30] ), .ZN(_00644_ ) );
AND2_X1 _07676_ ( .A1(_00644_ ), .A2(\u_idu.imm_auipc_lui [13] ), .ZN(_00645_ ) );
INV_X1 _07677_ ( .A(\u_idu.imm_auipc_lui [12] ), .ZN(_00646_ ) );
AND3_X1 _07678_ ( .A1(_00643_ ), .A2(_00645_ ), .A3(_00646_ ), .ZN(_00647_ ) );
INV_X1 _07679_ ( .A(\u_idu.imm_auipc_lui [14] ), .ZN(_00648_ ) );
NOR2_X1 _07680_ ( .A1(_00648_ ), .A2(\u_idu.imm_auipc_lui [25] ), .ZN(_00649_ ) );
NAND2_X1 _07681_ ( .A1(_00647_ ), .A2(_00649_ ), .ZN(_00650_ ) );
NOR2_X1 _07682_ ( .A1(\u_idu.imm_auipc_lui [14] ), .A2(\u_idu.imm_auipc_lui [25] ), .ZN(_00651_ ) );
NAND3_X1 _07683_ ( .A1(_00643_ ), .A2(_00645_ ), .A3(_00651_ ), .ZN(_00652_ ) );
AND2_X1 _07684_ ( .A1(_00650_ ), .A2(_00652_ ), .ZN(_00653_ ) );
AND3_X1 _07685_ ( .A1(_00641_ ), .A2(_00644_ ), .A3(_00642_ ), .ZN(_00654_ ) );
NOR2_X1 _07686_ ( .A1(\u_idu.imm_auipc_lui [12] ), .A2(\u_idu.imm_auipc_lui [13] ), .ZN(_00655_ ) );
INV_X1 _07687_ ( .A(\u_idu.imm_auipc_lui [25] ), .ZN(_00656_ ) );
AND3_X1 _07688_ ( .A1(_00655_ ), .A2(\u_idu.imm_auipc_lui [14] ), .A3(_00656_ ), .ZN(_00657_ ) );
NAND2_X1 _07689_ ( .A1(_00654_ ), .A2(_00657_ ), .ZN(_00658_ ) );
NAND4_X1 _07690_ ( .A1(_00643_ ), .A2(_00645_ ), .A3(\u_idu.imm_auipc_lui [12] ), .A4(_00649_ ), .ZN(_00659_ ) );
AND3_X1 _07691_ ( .A1(_00653_ ), .A2(_00658_ ), .A3(_00659_ ), .ZN(_00660_ ) );
AND3_X1 _07692_ ( .A1(_00643_ ), .A2(_00655_ ), .A3(_00651_ ), .ZN(_00661_ ) );
INV_X1 _07693_ ( .A(\u_idu.imm_auipc_lui [31] ), .ZN(_00662_ ) );
AND2_X1 _07694_ ( .A1(_00661_ ), .A2(_00662_ ), .ZN(_00663_ ) );
INV_X1 _07695_ ( .A(_00663_ ), .ZN(_00664_ ) );
NOR2_X1 _07696_ ( .A1(_00646_ ), .A2(\u_idu.imm_auipc_lui [13] ), .ZN(_00665_ ) );
AND3_X1 _07697_ ( .A1(_00654_ ), .A2(_00665_ ), .A3(_00651_ ), .ZN(_00666_ ) );
AND3_X1 _07698_ ( .A1(_00643_ ), .A2(_00665_ ), .A3(_00649_ ), .ZN(_00667_ ) );
AOI21_X1 _07699_ ( .A(_00666_ ), .B1(_00662_ ), .B2(_00667_ ), .ZN(_00668_ ) );
NAND3_X1 _07700_ ( .A1(_00660_ ), .A2(_00664_ ), .A3(_00668_ ), .ZN(_00669_ ) );
AND2_X4 _07701_ ( .A1(\u_idu.inst [0] ), .A2(\u_idu.inst [1] ), .ZN(_00670_ ) );
NOR2_X1 _07702_ ( .A1(\u_idu.inst [3] ), .A2(\u_idu.inst [2] ), .ZN(_00671_ ) );
AND2_X2 _07703_ ( .A1(_00670_ ), .A2(_00671_ ), .ZN(_00672_ ) );
INV_X1 _07704_ ( .A(\u_idu.inst [6] ), .ZN(_00673_ ) );
AND3_X1 _07705_ ( .A1(_00673_ ), .A2(\u_idu.inst [5] ), .A3(\u_idu.inst [4] ), .ZN(_00674_ ) );
AND2_X1 _07706_ ( .A1(_00672_ ), .A2(_00674_ ), .ZN(_00675_ ) );
AND2_X1 _07707_ ( .A1(_00669_ ), .A2(_00675_ ), .ZN(_00676_ ) );
NOR3_X1 _07708_ ( .A1(\u_idu.inst [5] ), .A2(\u_idu.inst [6] ), .A3(\u_idu.inst [4] ), .ZN(_00677_ ) );
AND2_X1 _07709_ ( .A1(_00672_ ), .A2(_00677_ ), .ZN(_00678_ ) );
OAI21_X1 _07710_ ( .A(\u_idu.imm_auipc_lui [13] ), .B1(\u_idu.imm_auipc_lui [12] ), .B2(\u_idu.imm_auipc_lui [14] ), .ZN(_00679_ ) );
AND2_X1 _07711_ ( .A1(_00678_ ), .A2(_00679_ ), .ZN(_00680_ ) );
NOR2_X1 _07712_ ( .A1(_00676_ ), .A2(_00680_ ), .ZN(_00681_ ) );
INV_X1 _07713_ ( .A(\u_idu.inst [5] ), .ZN(_00682_ ) );
NOR3_X1 _07714_ ( .A1(_00682_ ), .A2(\u_idu.inst [4] ), .A3(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ), .ZN(_00683_ ) );
AND2_X2 _07715_ ( .A1(_00672_ ), .A2(_00683_ ), .ZN(_00684_ ) );
NOR3_X1 _07716_ ( .A1(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A2(\u_idu.imm_auipc_lui [14] ), .A3(\u_idu.imm_auipc_lui [13] ), .ZN(_00685_ ) );
AOI21_X1 _07717_ ( .A(_00685_ ), .B1(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(\u_idu.imm_auipc_lui [13] ), .ZN(_00686_ ) );
AND2_X1 _07718_ ( .A1(_00684_ ), .A2(_00686_ ), .ZN(_00687_ ) );
INV_X1 _07719_ ( .A(_00687_ ), .ZN(_00688_ ) );
AND3_X1 _07720_ ( .A1(_00670_ ), .A2(_00673_ ), .A3(_00671_ ), .ZN(_00689_ ) );
INV_X1 _07721_ ( .A(\u_idu.inst [4] ), .ZN(_00690_ ) );
AND2_X1 _07722_ ( .A1(_00689_ ), .A2(_00690_ ), .ZN(_00691_ ) );
AND2_X1 _07723_ ( .A1(_00691_ ), .A2(\u_idu.inst [5] ), .ZN(_00692_ ) );
AND2_X2 _07724_ ( .A1(_00665_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00693_ ) );
INV_X1 _07725_ ( .A(_00693_ ), .ZN(_00694_ ) );
INV_X1 _07726_ ( .A(\u_idu.imm_auipc_lui [13] ), .ZN(_00695_ ) );
NOR2_X1 _07727_ ( .A1(_00695_ ), .A2(\u_idu.imm_auipc_lui [12] ), .ZN(_00696_ ) );
AND2_X1 _07728_ ( .A1(_00696_ ), .A2(_00648_ ), .ZN(_00697_ ) );
INV_X1 _07729_ ( .A(_00697_ ), .ZN(_00698_ ) );
AND2_X1 _07730_ ( .A1(_00655_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00699_ ) );
INV_X1 _07731_ ( .A(_00699_ ), .ZN(_00700_ ) );
NAND3_X1 _07732_ ( .A1(_00694_ ), .A2(_00698_ ), .A3(_00700_ ), .ZN(_00701_ ) );
AND2_X1 _07733_ ( .A1(_00692_ ), .A2(_00701_ ), .ZN(_00702_ ) );
NOR3_X1 _07734_ ( .A1(_00682_ ), .A2(_00690_ ), .A3(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ), .ZN(_00703_ ) );
AND2_X2 _07735_ ( .A1(_00672_ ), .A2(_00703_ ), .ZN(_00704_ ) );
INV_X1 _07736_ ( .A(_00704_ ), .ZN(_00705_ ) );
NOR2_X1 _07737_ ( .A1(_00693_ ), .A2(_00697_ ), .ZN(_00706_ ) );
NOR2_X1 _07738_ ( .A1(_00705_ ), .A2(_00706_ ), .ZN(_00707_ ) );
NOR2_X1 _07739_ ( .A1(_00702_ ), .A2(_00707_ ), .ZN(_00708_ ) );
AND3_X2 _07740_ ( .A1(_00681_ ), .A2(_00688_ ), .A3(_00708_ ), .ZN(_00709_ ) );
NOR3_X1 _07741_ ( .A1(_00690_ ), .A2(\u_idu.inst [5] ), .A3(\u_idu.inst [6] ), .ZN(_00710_ ) );
AND2_X2 _07742_ ( .A1(_00672_ ), .A2(_00710_ ), .ZN(_00711_ ) );
NAND3_X1 _07743_ ( .A1(\u_idu.inst [2] ), .A2(\u_idu.inst [0] ), .A3(\u_idu.inst [1] ), .ZN(_00712_ ) );
NOR2_X2 _07744_ ( .A1(_00712_ ), .A2(\u_idu.inst [3] ), .ZN(_00713_ ) );
NOR2_X1 _07745_ ( .A1(_00690_ ), .A2(\u_idu.inst [6] ), .ZN(_00714_ ) );
AND2_X1 _07746_ ( .A1(_00713_ ), .A2(_00714_ ), .ZN(_00715_ ) );
NOR2_X1 _07747_ ( .A1(_00711_ ), .A2(_00715_ ), .ZN(_00716_ ) );
AND2_X1 _07748_ ( .A1(_00713_ ), .A2(_00683_ ), .ZN(_00717_ ) );
BUF_X2 _07749_ ( .A(_00699_ ), .Z(_00718_ ) );
AND2_X2 _07750_ ( .A1(_00717_ ), .A2(_00718_ ), .ZN(_00719_ ) );
AND3_X1 _07751_ ( .A1(_00670_ ), .A2(\u_idu.inst [3] ), .A3(\u_idu.inst [2] ), .ZN(_00720_ ) );
AND2_X1 _07752_ ( .A1(_00720_ ), .A2(_00683_ ), .ZN(_00721_ ) );
NOR3_X1 _07753_ ( .A1(_00707_ ), .A2(_00719_ ), .A3(_00721_ ), .ZN(_00722_ ) );
AND3_X1 _07754_ ( .A1(_00681_ ), .A2(_00716_ ), .A3(_00722_ ), .ZN(_00723_ ) );
AND2_X1 _07755_ ( .A1(_00720_ ), .A2(_00677_ ), .ZN(_00724_ ) );
AND2_X1 _07756_ ( .A1(_00724_ ), .A2(_00694_ ), .ZN(_00725_ ) );
INV_X1 _07757_ ( .A(_00725_ ), .ZN(_00726_ ) );
AOI21_X1 _07758_ ( .A(_00711_ ), .B1(_00717_ ), .B2(_00718_ ), .ZN(_00727_ ) );
AND2_X1 _07759_ ( .A1(_00641_ ), .A2(_00644_ ), .ZN(_00728_ ) );
NOR2_X1 _07760_ ( .A1(\u_idu.imm_auipc_lui [22] ), .A2(fanout_net_20 ), .ZN(_00729_ ) );
AND2_X1 _07761_ ( .A1(_00728_ ), .A2(_00729_ ), .ZN(_00730_ ) );
NOR3_X4 _07762_ ( .A1(\u_idu.imm_auipc_lui [25] ), .A2(\u_idu.imm_auipc_lui [24] ), .A3(\u_idu.imm_auipc_lui [27] ), .ZN(_00731_ ) );
INV_X1 _07763_ ( .A(\u_idu.imm_auipc_lui [26] ), .ZN(_00732_ ) );
AND2_X1 _07764_ ( .A1(_00731_ ), .A2(_00732_ ), .ZN(_00733_ ) );
INV_X1 _07765_ ( .A(\u_idu.imm_auipc_lui [23] ), .ZN(_00734_ ) );
AND4_X1 _07766_ ( .A1(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A2(_00655_ ), .A3(_00734_ ), .A4(\u_idu.imm_auipc_lui [20] ), .ZN(_00735_ ) );
NAND4_X1 _07767_ ( .A1(_00704_ ), .A2(_00730_ ), .A3(_00733_ ), .A4(_00735_ ), .ZN(_00736_ ) );
AND3_X1 _07768_ ( .A1(_00726_ ), .A2(_00727_ ), .A3(_00736_ ), .ZN(_00737_ ) );
NAND3_X1 _07769_ ( .A1(_00709_ ), .A2(_00723_ ), .A3(_00737_ ), .ZN(_00738_ ) );
AND2_X1 _07770_ ( .A1(_00724_ ), .A2(_00693_ ), .ZN(_00739_ ) );
AOI211_X1 _07771_ ( .A(_00680_ ), .B(_00739_ ), .C1(_00669_ ), .C2(_00675_ ), .ZN(_00740_ ) );
AOI211_X1 _07772_ ( .A(_00719_ ), .B(_00707_ ), .C1(_00692_ ), .C2(_00701_ ), .ZN(_00741_ ) );
AND3_X1 _07773_ ( .A1(_00740_ ), .A2(_00716_ ), .A3(_00741_ ), .ZN(_00742_ ) );
NOR2_X1 _07774_ ( .A1(_00719_ ), .A2(_00721_ ), .ZN(_00743_ ) );
INV_X1 _07775_ ( .A(_00743_ ), .ZN(_00744_ ) );
OR2_X1 _07776_ ( .A1(_00742_ ), .A2(_00744_ ), .ZN(_00745_ ) );
NAND2_X1 _07777_ ( .A1(_00738_ ), .A2(_00745_ ), .ZN(_00746_ ) );
AND2_X1 _07778_ ( .A1(_00704_ ), .A2(_00718_ ), .ZN(_00747_ ) );
INV_X1 _07779_ ( .A(\u_idu.imm_auipc_lui [20] ), .ZN(_00748_ ) );
BUF_X2 _07780_ ( .A(_00748_ ), .Z(_00749_ ) );
AND3_X1 _07781_ ( .A1(_00731_ ), .A2(_00734_ ), .A3(_00732_ ), .ZN(_00750_ ) );
AND3_X1 _07782_ ( .A1(_00747_ ), .A2(_00749_ ), .A3(_00750_ ), .ZN(_00751_ ) );
AND2_X1 _07783_ ( .A1(\u_idu.imm_auipc_lui [28] ), .A2(\u_idu.imm_auipc_lui [29] ), .ZN(_00752_ ) );
AND2_X1 _07784_ ( .A1(_00752_ ), .A2(_00644_ ), .ZN(_00753_ ) );
BUF_X4 _07785_ ( .A(_00753_ ), .Z(_00754_ ) );
INV_X1 _07786_ ( .A(fanout_net_20 ), .ZN(_00755_ ) );
NOR2_X1 _07787_ ( .A1(_00755_ ), .A2(\u_idu.imm_auipc_lui [22] ), .ZN(_00756_ ) );
AND2_X1 _07788_ ( .A1(_00754_ ), .A2(_00756_ ), .ZN(_00757_ ) );
AOI21_X1 _07789_ ( .A(_00739_ ), .B1(_00751_ ), .B2(_00757_ ), .ZN(_00758_ ) );
AND2_X1 _07790_ ( .A1(_00746_ ), .A2(_00758_ ), .ZN(_00759_ ) );
CLKBUF_X2 _07791_ ( .A(_00637_ ), .Z(_00760_ ) );
INV_X1 _07792_ ( .A(_00760_ ), .ZN(_00761_ ) );
INV_X1 _07793_ ( .A(\u_exu.eopt [12] ), .ZN(_00762_ ) );
OR4_X1 _07794_ ( .A1(\ea_mask [1] ), .A2(_00762_ ), .A3(\ea_mask [0] ), .A4(\u_exu.eopt [15] ), .ZN(_00763_ ) );
NOR3_X2 _07795_ ( .A1(_00761_ ), .A2(\u_exu.eopt [0] ), .A3(_00763_ ), .ZN(_00764_ ) );
NOR2_X1 _07796_ ( .A1(_00764_ ), .A2(\u_exu.jmpc_ok ), .ZN(_00765_ ) );
OAI21_X1 _07797_ ( .A(_00640_ ), .B1(_00759_ ), .B2(_00765_ ), .ZN(_00766_ ) );
INV_X1 _07798_ ( .A(exe_valid ), .ZN(_00767_ ) );
AND2_X1 _07799_ ( .A1(_00767_ ), .A2(idu_ready ), .ZN(_00768_ ) );
BUF_X4 _07800_ ( .A(_00768_ ), .Z(_00769_ ) );
BUF_X4 _07801_ ( .A(_00769_ ), .Z(_00770_ ) );
OR2_X1 _07802_ ( .A1(_00766_ ), .A2(_00770_ ), .ZN(_00000_ ) );
INV_X1 _07803_ ( .A(fanout_net_1 ), .ZN(_00771_ ) );
BUF_X2 _07804_ ( .A(_00771_ ), .Z(_00772_ ) );
CLKBUF_X2 _07805_ ( .A(_00772_ ), .Z(_00773_ ) );
AND2_X1 _07806_ ( .A1(_00773_ ), .A2(\ea_addr [31] ), .ZN(_00001_ ) );
AND2_X1 _07807_ ( .A1(_00773_ ), .A2(\ea_addr [30] ), .ZN(_00002_ ) );
AND2_X1 _07808_ ( .A1(_00773_ ), .A2(\ea_addr [21] ), .ZN(_00003_ ) );
AND2_X1 _07809_ ( .A1(_00773_ ), .A2(\ea_addr [20] ), .ZN(_00004_ ) );
AND2_X1 _07810_ ( .A1(_00773_ ), .A2(\ea_addr [19] ), .ZN(_00005_ ) );
AND2_X1 _07811_ ( .A1(_00773_ ), .A2(\ea_addr [18] ), .ZN(_00006_ ) );
AND2_X1 _07812_ ( .A1(_00773_ ), .A2(\ea_addr [17] ), .ZN(_00007_ ) );
CLKBUF_X2 _07813_ ( .A(_00772_ ), .Z(_00774_ ) );
AND2_X1 _07814_ ( .A1(_00774_ ), .A2(\ea_addr [16] ), .ZN(_00008_ ) );
AND2_X1 _07815_ ( .A1(_00774_ ), .A2(\ea_addr [15] ), .ZN(_00009_ ) );
AND2_X1 _07816_ ( .A1(_00774_ ), .A2(\ea_addr [14] ), .ZN(_00010_ ) );
AND2_X1 _07817_ ( .A1(_00774_ ), .A2(\ea_addr [13] ), .ZN(_00011_ ) );
AND2_X1 _07818_ ( .A1(_00774_ ), .A2(\ea_addr [12] ), .ZN(_00012_ ) );
AND2_X1 _07819_ ( .A1(_00774_ ), .A2(\ea_addr [29] ), .ZN(_00013_ ) );
AND2_X1 _07820_ ( .A1(_00774_ ), .A2(\ea_addr [11] ), .ZN(_00014_ ) );
AND2_X1 _07821_ ( .A1(_00774_ ), .A2(\ea_addr [10] ), .ZN(_00015_ ) );
AND2_X1 _07822_ ( .A1(_00774_ ), .A2(\ea_addr [9] ), .ZN(_00016_ ) );
AND2_X1 _07823_ ( .A1(_00774_ ), .A2(\ea_addr [8] ), .ZN(_00017_ ) );
CLKBUF_X2 _07824_ ( .A(_00772_ ), .Z(_00775_ ) );
AND2_X1 _07825_ ( .A1(_00775_ ), .A2(\ea_addr [7] ), .ZN(_00018_ ) );
AND2_X1 _07826_ ( .A1(_00775_ ), .A2(\ea_addr [6] ), .ZN(_00019_ ) );
AND2_X1 _07827_ ( .A1(_00775_ ), .A2(\ea_addr [5] ), .ZN(_00020_ ) );
AND2_X1 _07828_ ( .A1(_00775_ ), .A2(\ea_addr [4] ), .ZN(_00021_ ) );
AND2_X1 _07829_ ( .A1(_00775_ ), .A2(\ea_addr [3] ), .ZN(_00022_ ) );
AND2_X1 _07830_ ( .A1(_00775_ ), .A2(\ea_addr [2] ), .ZN(_00023_ ) );
AND2_X1 _07831_ ( .A1(_00775_ ), .A2(\ea_addr [28] ), .ZN(_00024_ ) );
AND2_X1 _07832_ ( .A1(_00775_ ), .A2(\ea_addr [1] ), .ZN(_00025_ ) );
AND2_X1 _07833_ ( .A1(_00775_ ), .A2(\ea_addr [0] ), .ZN(_00026_ ) );
AND2_X1 _07834_ ( .A1(_00775_ ), .A2(\ea_addr [27] ), .ZN(_00027_ ) );
CLKBUF_X2 _07835_ ( .A(_00772_ ), .Z(_00776_ ) );
AND2_X1 _07836_ ( .A1(_00776_ ), .A2(\ea_addr [26] ), .ZN(_00028_ ) );
AND2_X1 _07837_ ( .A1(_00776_ ), .A2(\ea_addr [25] ), .ZN(_00029_ ) );
AND2_X1 _07838_ ( .A1(_00776_ ), .A2(\ea_addr [24] ), .ZN(_00030_ ) );
AND2_X1 _07839_ ( .A1(_00776_ ), .A2(\ea_addr [23] ), .ZN(_00031_ ) );
AND2_X1 _07840_ ( .A1(_00776_ ), .A2(\ea_addr [22] ), .ZN(_00032_ ) );
NOR2_X1 _07841_ ( .A1(_00629_ ), .A2(fanout_net_1 ), .ZN(_00033_ ) );
NOR2_X1 _07842_ ( .A1(_00630_ ), .A2(fanout_net_1 ), .ZN(_00034_ ) );
AND2_X1 _07843_ ( .A1(_00776_ ), .A2(ea_rsign ), .ZN(_00035_ ) );
AND2_X1 _07844_ ( .A1(_00631_ ), .A2(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ), .ZN(_00777_ ) );
AND3_X1 _07845_ ( .A1(_00760_ ), .A2(\u_exu.eopt [12] ), .A3(_00777_ ), .ZN(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_AND__A_Y ) );
CLKBUF_X2 _07846_ ( .A(_00771_ ), .Z(_00778_ ) );
AND4_X1 _07847_ ( .A1(_00778_ ), .A2(_00760_ ), .A3(\u_exu.eopt [12] ), .A4(_00777_ ), .ZN(_00036_ ) );
AND2_X1 _07848_ ( .A1(_00776_ ), .A2(\ea_ard [3] ), .ZN(_00037_ ) );
AND2_X1 _07849_ ( .A1(_00776_ ), .A2(\ea_ard [2] ), .ZN(_00038_ ) );
AND2_X1 _07850_ ( .A1(_00776_ ), .A2(\ea_ard [1] ), .ZN(_00039_ ) );
AND2_X1 _07851_ ( .A1(_00776_ ), .A2(\ea_ard [0] ), .ZN(_00040_ ) );
CLKBUF_X2 _07852_ ( .A(_00772_ ), .Z(_00779_ ) );
AND2_X1 _07853_ ( .A1(_00779_ ), .A2(\ea_wdata [31] ), .ZN(_00041_ ) );
AND2_X1 _07854_ ( .A1(_00779_ ), .A2(\ea_wdata [30] ), .ZN(_00042_ ) );
AND2_X1 _07855_ ( .A1(_00779_ ), .A2(\ea_wdata [21] ), .ZN(_00043_ ) );
AND2_X1 _07856_ ( .A1(_00779_ ), .A2(\ea_wdata [20] ), .ZN(_00044_ ) );
AND2_X1 _07857_ ( .A1(_00779_ ), .A2(\ea_wdata [19] ), .ZN(_00045_ ) );
AND2_X1 _07858_ ( .A1(_00779_ ), .A2(\ea_wdata [18] ), .ZN(_00046_ ) );
AND2_X1 _07859_ ( .A1(_00779_ ), .A2(\ea_wdata [17] ), .ZN(_00047_ ) );
AND2_X1 _07860_ ( .A1(_00779_ ), .A2(\ea_wdata [16] ), .ZN(_00048_ ) );
AND2_X1 _07861_ ( .A1(_00779_ ), .A2(\ea_wdata [15] ), .ZN(_00049_ ) );
AND2_X1 _07862_ ( .A1(_00779_ ), .A2(\ea_wdata [14] ), .ZN(_00050_ ) );
CLKBUF_X2 _07863_ ( .A(_00772_ ), .Z(_00780_ ) );
AND2_X1 _07864_ ( .A1(_00780_ ), .A2(\ea_wdata [13] ), .ZN(_00051_ ) );
AND2_X1 _07865_ ( .A1(_00780_ ), .A2(\ea_wdata [12] ), .ZN(_00052_ ) );
AND2_X1 _07866_ ( .A1(_00780_ ), .A2(\ea_wdata [29] ), .ZN(_00053_ ) );
AND2_X1 _07867_ ( .A1(_00780_ ), .A2(\ea_wdata [11] ), .ZN(_00054_ ) );
AND2_X1 _07868_ ( .A1(_00780_ ), .A2(\ea_wdata [10] ), .ZN(_00055_ ) );
AND2_X1 _07869_ ( .A1(_00780_ ), .A2(\ea_wdata [9] ), .ZN(_00056_ ) );
AND2_X1 _07870_ ( .A1(_00780_ ), .A2(\ea_wdata [8] ), .ZN(_00057_ ) );
AND2_X1 _07871_ ( .A1(_00780_ ), .A2(\ea_wdata [7] ), .ZN(_00058_ ) );
AND2_X1 _07872_ ( .A1(_00780_ ), .A2(\ea_wdata [6] ), .ZN(_00059_ ) );
AND2_X1 _07873_ ( .A1(_00780_ ), .A2(\ea_wdata [5] ), .ZN(_00060_ ) );
CLKBUF_X2 _07874_ ( .A(_00772_ ), .Z(_00781_ ) );
AND2_X1 _07875_ ( .A1(_00781_ ), .A2(\ea_wdata [4] ), .ZN(_00061_ ) );
AND2_X1 _07876_ ( .A1(_00781_ ), .A2(\ea_wdata [3] ), .ZN(_00062_ ) );
AND2_X1 _07877_ ( .A1(_00781_ ), .A2(\ea_wdata [2] ), .ZN(_00063_ ) );
AND2_X1 _07878_ ( .A1(_00781_ ), .A2(\ea_wdata [28] ), .ZN(_00064_ ) );
AND2_X1 _07879_ ( .A1(_00781_ ), .A2(\ea_wdata [1] ), .ZN(_00065_ ) );
AND2_X1 _07880_ ( .A1(_00781_ ), .A2(\ea_wdata [0] ), .ZN(_00066_ ) );
AND2_X1 _07881_ ( .A1(_00781_ ), .A2(\ea_wdata [27] ), .ZN(_00067_ ) );
AND2_X1 _07882_ ( .A1(_00781_ ), .A2(\ea_wdata [26] ), .ZN(_00068_ ) );
AND2_X1 _07883_ ( .A1(_00781_ ), .A2(\ea_wdata [25] ), .ZN(_00069_ ) );
AND2_X1 _07884_ ( .A1(_00781_ ), .A2(\ea_wdata [24] ), .ZN(_00070_ ) );
CLKBUF_X2 _07885_ ( .A(_00771_ ), .Z(_00782_ ) );
AND2_X1 _07886_ ( .A1(_00782_ ), .A2(\ea_wdata [23] ), .ZN(_00071_ ) );
AND2_X1 _07887_ ( .A1(_00782_ ), .A2(\ea_wdata [22] ), .ZN(_00072_ ) );
INV_X1 _07888_ ( .A(_00777_ ), .ZN(_00783_ ) );
NOR4_X1 _07889_ ( .A1(_00633_ ), .A2(fanout_net_1 ), .A3(_00636_ ), .A4(_00783_ ), .ZN(_00073_ ) );
AND3_X1 _07890_ ( .A1(_00760_ ), .A2(_00762_ ), .A3(_00777_ ), .ZN(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND4_X1 _07891_ ( .A1(_00778_ ), .A2(_00760_ ), .A3(_00762_ ), .A4(_00777_ ), .ZN(_00074_ ) );
INV_X1 _07892_ ( .A(fanout_net_5 ), .ZN(_00784_ ) );
BUF_X2 _07893_ ( .A(_00784_ ), .Z(_00785_ ) );
OR2_X1 _07894_ ( .A1(_00785_ ), .A2(\ea_pc [31] ), .ZN(_00786_ ) );
OR2_X1 _07895_ ( .A1(\ea_addr [31] ), .A2(fanout_net_5 ), .ZN(_00787_ ) );
AND3_X1 _07896_ ( .A1(_00786_ ), .A2(_00782_ ), .A3(_00787_ ), .ZN(_00075_ ) );
CLKBUF_X2 _07897_ ( .A(_00785_ ), .Z(_00788_ ) );
BUF_X2 _07898_ ( .A(_00788_ ), .Z(_00789_ ) );
OR2_X1 _07899_ ( .A1(_00789_ ), .A2(\ea_pc [30] ), .ZN(_00790_ ) );
OR2_X1 _07900_ ( .A1(\ea_addr [30] ), .A2(fanout_net_5 ), .ZN(_00791_ ) );
AND3_X1 _07901_ ( .A1(_00790_ ), .A2(_00782_ ), .A3(_00791_ ), .ZN(_00076_ ) );
OR2_X1 _07902_ ( .A1(_00785_ ), .A2(\ea_pc [21] ), .ZN(_00792_ ) );
OR2_X1 _07903_ ( .A1(\ea_addr [21] ), .A2(fanout_net_5 ), .ZN(_00793_ ) );
AND3_X1 _07904_ ( .A1(_00792_ ), .A2(_00782_ ), .A3(_00793_ ), .ZN(_00077_ ) );
OR2_X1 _07905_ ( .A1(_00788_ ), .A2(\ea_pc [20] ), .ZN(_00794_ ) );
OR2_X1 _07906_ ( .A1(\ea_addr [20] ), .A2(fanout_net_5 ), .ZN(_00795_ ) );
AND3_X1 _07907_ ( .A1(_00794_ ), .A2(_00782_ ), .A3(_00795_ ), .ZN(_00078_ ) );
OR2_X1 _07908_ ( .A1(_00788_ ), .A2(\ea_pc [19] ), .ZN(_00796_ ) );
OR2_X1 _07909_ ( .A1(\ea_addr [19] ), .A2(fanout_net_5 ), .ZN(_00797_ ) );
AND3_X1 _07910_ ( .A1(_00796_ ), .A2(_00782_ ), .A3(_00797_ ), .ZN(_00079_ ) );
CLKBUF_X2 _07911_ ( .A(_00785_ ), .Z(_00798_ ) );
OR2_X1 _07912_ ( .A1(_00798_ ), .A2(\ea_pc [18] ), .ZN(_00799_ ) );
OR2_X1 _07913_ ( .A1(\ea_addr [18] ), .A2(fanout_net_5 ), .ZN(_00800_ ) );
AND3_X1 _07914_ ( .A1(_00799_ ), .A2(_00782_ ), .A3(_00800_ ), .ZN(_00080_ ) );
OR2_X1 _07915_ ( .A1(_00788_ ), .A2(\ea_pc [17] ), .ZN(_00801_ ) );
OR2_X1 _07916_ ( .A1(\ea_addr [17] ), .A2(fanout_net_5 ), .ZN(_00802_ ) );
AND3_X1 _07917_ ( .A1(_00801_ ), .A2(_00782_ ), .A3(_00802_ ), .ZN(_00081_ ) );
OR2_X1 _07918_ ( .A1(_00788_ ), .A2(\ea_pc [16] ), .ZN(_00803_ ) );
OR2_X1 _07919_ ( .A1(\ea_addr [16] ), .A2(fanout_net_5 ), .ZN(_00804_ ) );
AND3_X1 _07920_ ( .A1(_00803_ ), .A2(_00782_ ), .A3(_00804_ ), .ZN(_00082_ ) );
OR2_X1 _07921_ ( .A1(_00798_ ), .A2(\ea_pc [15] ), .ZN(_00805_ ) );
CLKBUF_X2 _07922_ ( .A(_00771_ ), .Z(_00806_ ) );
OR2_X1 _07923_ ( .A1(\ea_addr [15] ), .A2(fanout_net_5 ), .ZN(_00807_ ) );
AND3_X1 _07924_ ( .A1(_00805_ ), .A2(_00806_ ), .A3(_00807_ ), .ZN(_00083_ ) );
OR2_X1 _07925_ ( .A1(_00788_ ), .A2(\ea_pc [14] ), .ZN(_00808_ ) );
OR2_X1 _07926_ ( .A1(\ea_addr [14] ), .A2(fanout_net_5 ), .ZN(_00809_ ) );
AND3_X1 _07927_ ( .A1(_00808_ ), .A2(_00806_ ), .A3(_00809_ ), .ZN(_00084_ ) );
OR2_X1 _07928_ ( .A1(_00798_ ), .A2(\ea_pc [13] ), .ZN(_00810_ ) );
OR2_X1 _07929_ ( .A1(\ea_addr [13] ), .A2(fanout_net_5 ), .ZN(_00811_ ) );
AND3_X1 _07930_ ( .A1(_00810_ ), .A2(_00806_ ), .A3(_00811_ ), .ZN(_00085_ ) );
OR2_X1 _07931_ ( .A1(_00798_ ), .A2(\ea_pc [10] ), .ZN(_00812_ ) );
OR2_X1 _07932_ ( .A1(\ea_addr [10] ), .A2(fanout_net_5 ), .ZN(_00813_ ) );
AND3_X1 _07933_ ( .A1(_00812_ ), .A2(_00806_ ), .A3(_00813_ ), .ZN(_00086_ ) );
OR2_X1 _07934_ ( .A1(_00798_ ), .A2(\ea_pc [29] ), .ZN(_00814_ ) );
OR2_X1 _07935_ ( .A1(\ea_addr [29] ), .A2(fanout_net_5 ), .ZN(_00815_ ) );
AND3_X1 _07936_ ( .A1(_00814_ ), .A2(_00806_ ), .A3(_00815_ ), .ZN(_00087_ ) );
OR2_X1 _07937_ ( .A1(_00798_ ), .A2(\ea_pc [9] ), .ZN(_00816_ ) );
OR2_X1 _07938_ ( .A1(\ea_addr [9] ), .A2(fanout_net_5 ), .ZN(_00817_ ) );
AND3_X1 _07939_ ( .A1(_00816_ ), .A2(_00806_ ), .A3(_00817_ ), .ZN(_00088_ ) );
OR2_X1 _07940_ ( .A1(_00788_ ), .A2(\ea_pc [8] ), .ZN(_00818_ ) );
OR2_X1 _07941_ ( .A1(\ea_addr [8] ), .A2(fanout_net_5 ), .ZN(_00819_ ) );
AND3_X1 _07942_ ( .A1(_00818_ ), .A2(_00806_ ), .A3(_00819_ ), .ZN(_00089_ ) );
OR2_X1 _07943_ ( .A1(_00788_ ), .A2(\ea_pc [7] ), .ZN(_00820_ ) );
OR2_X1 _07944_ ( .A1(\ea_addr [7] ), .A2(fanout_net_5 ), .ZN(_00821_ ) );
AND3_X1 _07945_ ( .A1(_00820_ ), .A2(_00806_ ), .A3(_00821_ ), .ZN(_00090_ ) );
OR2_X1 _07946_ ( .A1(_00798_ ), .A2(\ea_pc [6] ), .ZN(_00822_ ) );
OR2_X1 _07947_ ( .A1(\ea_addr [6] ), .A2(fanout_net_5 ), .ZN(_00823_ ) );
AND3_X1 _07948_ ( .A1(_00822_ ), .A2(_00806_ ), .A3(_00823_ ), .ZN(_00091_ ) );
NAND2_X1 _07949_ ( .A1(_00789_ ), .A2(\ea_addr [5] ), .ZN(_00824_ ) );
NAND2_X1 _07950_ ( .A1(fanout_net_5 ), .A2(\ea_pc [5] ), .ZN(_00825_ ) );
AOI21_X1 _07951_ ( .A(fanout_net_1 ), .B1(_00824_ ), .B2(_00825_ ), .ZN(_00092_ ) );
OR2_X1 _07952_ ( .A1(_00789_ ), .A2(\ea_pc [4] ), .ZN(_00826_ ) );
OR2_X1 _07953_ ( .A1(\ea_addr [4] ), .A2(fanout_net_5 ), .ZN(_00827_ ) );
AND3_X1 _07954_ ( .A1(_00826_ ), .A2(_00806_ ), .A3(_00827_ ), .ZN(_00093_ ) );
OR2_X1 _07955_ ( .A1(_00798_ ), .A2(\ea_pc [3] ), .ZN(_00828_ ) );
CLKBUF_X2 _07956_ ( .A(_00771_ ), .Z(_00829_ ) );
OR2_X1 _07957_ ( .A1(\ea_addr [3] ), .A2(fanout_net_5 ), .ZN(_00830_ ) );
AND3_X1 _07958_ ( .A1(_00828_ ), .A2(_00829_ ), .A3(_00830_ ), .ZN(_00094_ ) );
NAND2_X1 _07959_ ( .A1(_00788_ ), .A2(\ea_addr [2] ), .ZN(_00831_ ) );
NAND2_X1 _07960_ ( .A1(fanout_net_5 ), .A2(\ea_pc [2] ), .ZN(_00832_ ) );
AOI21_X1 _07961_ ( .A(fanout_net_1 ), .B1(_00831_ ), .B2(_00832_ ), .ZN(_00095_ ) );
NAND2_X1 _07962_ ( .A1(_00789_ ), .A2(\ea_addr [1] ), .ZN(_00833_ ) );
NAND2_X1 _07963_ ( .A1(fanout_net_5 ), .A2(\ea_pc [1] ), .ZN(_00834_ ) );
AOI21_X1 _07964_ ( .A(fanout_net_1 ), .B1(_00833_ ), .B2(_00834_ ), .ZN(_00096_ ) );
NAND2_X1 _07965_ ( .A1(_00785_ ), .A2(\ea_addr [0] ), .ZN(_00835_ ) );
NAND2_X1 _07966_ ( .A1(fanout_net_5 ), .A2(\ea_pc [0] ), .ZN(_00836_ ) );
AOI21_X1 _07967_ ( .A(fanout_net_1 ), .B1(_00835_ ), .B2(_00836_ ), .ZN(_00097_ ) );
OR2_X1 _07968_ ( .A1(_00789_ ), .A2(\ea_pc [28] ), .ZN(_00837_ ) );
OR2_X1 _07969_ ( .A1(\ea_addr [28] ), .A2(fanout_net_5 ), .ZN(_00838_ ) );
AND3_X1 _07970_ ( .A1(_00837_ ), .A2(_00829_ ), .A3(_00838_ ), .ZN(_00098_ ) );
OR2_X1 _07971_ ( .A1(_00798_ ), .A2(\ea_pc [27] ), .ZN(_00839_ ) );
OR2_X1 _07972_ ( .A1(\ea_addr [27] ), .A2(fanout_net_5 ), .ZN(_00840_ ) );
AND3_X1 _07973_ ( .A1(_00839_ ), .A2(_00829_ ), .A3(_00840_ ), .ZN(_00099_ ) );
NAND2_X1 _07974_ ( .A1(_00789_ ), .A2(\ea_addr [26] ), .ZN(_00841_ ) );
NAND2_X1 _07975_ ( .A1(fanout_net_5 ), .A2(\ea_pc [26] ), .ZN(_00842_ ) );
AOI21_X1 _07976_ ( .A(fanout_net_1 ), .B1(_00841_ ), .B2(_00842_ ), .ZN(_00100_ ) );
OR2_X1 _07977_ ( .A1(_00798_ ), .A2(\ea_pc [25] ), .ZN(_00843_ ) );
OR2_X1 _07978_ ( .A1(\ea_addr [25] ), .A2(fanout_net_5 ), .ZN(_00844_ ) );
AND3_X1 _07979_ ( .A1(_00843_ ), .A2(_00829_ ), .A3(_00844_ ), .ZN(_00101_ ) );
OR2_X1 _07980_ ( .A1(_00785_ ), .A2(\ea_pc [24] ), .ZN(_00845_ ) );
OR2_X1 _07981_ ( .A1(\ea_addr [24] ), .A2(ea_err ), .ZN(_00846_ ) );
AND3_X1 _07982_ ( .A1(_00845_ ), .A2(_00829_ ), .A3(_00846_ ), .ZN(_00102_ ) );
NAND2_X1 _07983_ ( .A1(_00789_ ), .A2(\ea_addr [23] ), .ZN(_00847_ ) );
NAND2_X1 _07984_ ( .A1(ea_err ), .A2(\ea_pc [23] ), .ZN(_00848_ ) );
AOI21_X1 _07985_ ( .A(fanout_net_1 ), .B1(_00847_ ), .B2(_00848_ ), .ZN(_00103_ ) );
OR2_X1 _07986_ ( .A1(_00785_ ), .A2(\ea_pc [22] ), .ZN(_00849_ ) );
OR2_X1 _07987_ ( .A1(\ea_addr [22] ), .A2(ea_err ), .ZN(_00850_ ) );
AND3_X1 _07988_ ( .A1(_00849_ ), .A2(_00829_ ), .A3(_00850_ ), .ZN(_00104_ ) );
NAND2_X1 _07989_ ( .A1(_00789_ ), .A2(\ea_addr [12] ), .ZN(_00851_ ) );
NAND2_X1 _07990_ ( .A1(ea_err ), .A2(\ea_pc [12] ), .ZN(_00852_ ) );
NAND3_X1 _07991_ ( .A1(_00851_ ), .A2(_00773_ ), .A3(_00852_ ), .ZN(_00105_ ) );
NAND2_X1 _07992_ ( .A1(_00789_ ), .A2(\ea_addr [11] ), .ZN(_00853_ ) );
NAND2_X1 _07993_ ( .A1(ea_err ), .A2(\ea_pc [11] ), .ZN(_00854_ ) );
NAND3_X1 _07994_ ( .A1(_00853_ ), .A2(_00773_ ), .A3(_00854_ ), .ZN(_00106_ ) );
AOI21_X1 _07995_ ( .A(fanout_net_1 ), .B1(_00851_ ), .B2(_00852_ ), .ZN(_00107_ ) );
AOI21_X1 _07996_ ( .A(fanout_net_1 ), .B1(_00853_ ), .B2(_00854_ ), .ZN(_00108_ ) );
BUF_X8 _07997_ ( .A(_00764_ ), .Z(_00855_ ) );
BUF_X4 _07998_ ( .A(_00855_ ), .Z(_00856_ ) );
BUF_X4 _07999_ ( .A(_00638_ ), .Z(_00857_ ) );
BUF_X4 _08000_ ( .A(_00857_ ), .Z(_00858_ ) );
BUF_X4 _08001_ ( .A(_00858_ ), .Z(_00859_ ) );
BUF_X2 _08002_ ( .A(_00662_ ), .Z(_00860_ ) );
NOR4_X1 _08003_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .A3(_00859_ ), .A4(_00860_ ), .ZN(_00110_ ) );
INV_X1 _08004_ ( .A(\u_idu.imm_auipc_lui [30] ), .ZN(_00861_ ) );
NOR4_X1 _08005_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .A3(_00859_ ), .A4(_00861_ ), .ZN(_00111_ ) );
NOR2_X1 _08006_ ( .A1(_00764_ ), .A2(fanout_net_1 ), .ZN(_00862_ ) );
BUF_X2 _08007_ ( .A(_00862_ ), .Z(_00863_ ) );
CLKBUF_X2 _08008_ ( .A(_00863_ ), .Z(_00864_ ) );
BUF_X2 _08009_ ( .A(_00640_ ), .Z(_00865_ ) );
CLKBUF_X2 _08010_ ( .A(_00865_ ), .Z(_00866_ ) );
AND3_X1 _08011_ ( .A1(_00655_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(\u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ), .ZN(_00867_ ) );
AND2_X2 _08012_ ( .A1(_00750_ ), .A2(_00867_ ), .ZN(_00868_ ) );
AND2_X1 _08013_ ( .A1(_00868_ ), .A2(_00757_ ), .ZN(_00869_ ) );
AND3_X1 _08014_ ( .A1(_00730_ ), .A2(_00733_ ), .A3(_00735_ ), .ZN(_00870_ ) );
NOR2_X2 _08015_ ( .A1(_00869_ ), .A2(_00870_ ), .ZN(_00871_ ) );
AND2_X1 _08016_ ( .A1(_00871_ ), .A2(fanout_net_20 ), .ZN(_00872_ ) );
AND3_X1 _08017_ ( .A1(_00864_ ), .A2(_00866_ ), .A3(_00872_ ), .ZN(_00112_ ) );
NAND3_X1 _08018_ ( .A1(_00757_ ), .A2(_00750_ ), .A3(_00867_ ), .ZN(_00873_ ) );
AND4_X1 _08019_ ( .A1(_00734_ ), .A2(_00731_ ), .A3(\u_idu.imm_auipc_lui [20] ), .A4(_00732_ ), .ZN(_00874_ ) );
NAND3_X1 _08020_ ( .A1(_00730_ ), .A2(_00718_ ), .A3(_00874_ ), .ZN(_00875_ ) );
AND2_X1 _08021_ ( .A1(_00873_ ), .A2(_00875_ ), .ZN(_00876_ ) );
NAND2_X1 _08022_ ( .A1(_00876_ ), .A2(\u_idu.imm_auipc_lui [20] ), .ZN(_00877_ ) );
NOR4_X1 _08023_ ( .A1(_00856_ ), .A2(_00877_ ), .A3(_00859_ ), .A4(fanout_net_1 ), .ZN(_00113_ ) );
NOR2_X1 _08024_ ( .A1(_00857_ ), .A2(fanout_net_1 ), .ZN(_00878_ ) );
INV_X1 _08025_ ( .A(_00878_ ), .ZN(_00879_ ) );
BUF_X4 _08026_ ( .A(_00879_ ), .Z(_00880_ ) );
BUF_X2 _08027_ ( .A(_00880_ ), .Z(flush_$_OR__Y_B ) );
INV_X1 _08028_ ( .A(\u_idu.imm_auipc_lui [29] ), .ZN(_00881_ ) );
BUF_X4 _08029_ ( .A(_00764_ ), .Z(_00882_ ) );
INV_X1 _08030_ ( .A(_00876_ ), .ZN(_00883_ ) );
NOR4_X1 _08031_ ( .A1(flush_$_OR__Y_B ), .A2(_00881_ ), .A3(_00882_ ), .A4(_00883_ ), .ZN(_00114_ ) );
INV_X1 _08032_ ( .A(\u_idu.imm_auipc_lui [28] ), .ZN(_00884_ ) );
NOR4_X1 _08033_ ( .A1(flush_$_OR__Y_B ), .A2(_00884_ ), .A3(_00882_ ), .A4(_00883_ ), .ZN(_00115_ ) );
BUF_X4 _08034_ ( .A(_00858_ ), .Z(_00885_ ) );
INV_X1 _08035_ ( .A(\u_idu.imm_auipc_lui [27] ), .ZN(_00886_ ) );
NOR4_X1 _08036_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_00886_ ), .ZN(_00116_ ) );
NOR4_X1 _08037_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_00732_ ), .ZN(_00117_ ) );
NOR4_X1 _08038_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_00656_ ), .ZN(_00118_ ) );
INV_X1 _08039_ ( .A(\u_idu.imm_auipc_lui [24] ), .ZN(_00887_ ) );
NOR4_X1 _08040_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_00887_ ), .ZN(_00119_ ) );
BUF_X2 _08041_ ( .A(_00734_ ), .Z(_00888_ ) );
NOR4_X1 _08042_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_00888_ ), .ZN(_00120_ ) );
BUF_X4 _08043_ ( .A(_00855_ ), .Z(_00889_ ) );
INV_X2 _08044_ ( .A(\u_idu.imm_auipc_lui [22] ), .ZN(_00890_ ) );
NOR4_X1 _08045_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_00890_ ), .ZN(_00121_ ) );
NOR2_X1 _08046_ ( .A1(_00879_ ), .A2(_00764_ ), .ZN(_00891_ ) );
INV_X1 _08047_ ( .A(_00891_ ), .ZN(_00892_ ) );
BUF_X4 _08048_ ( .A(_00892_ ), .Z(_00893_ ) );
BUF_X4 _08049_ ( .A(_00893_ ), .Z(_00894_ ) );
NOR2_X2 _08050_ ( .A1(_00721_ ), .A2(_00678_ ), .ZN(_00895_ ) );
INV_X1 _08051_ ( .A(_00675_ ), .ZN(_00896_ ) );
NAND3_X1 _08052_ ( .A1(_00895_ ), .A2(_00705_ ), .A3(_00896_ ), .ZN(_00897_ ) );
INV_X2 _08053_ ( .A(_00711_ ), .ZN(_00898_ ) );
INV_X1 _08054_ ( .A(_00717_ ), .ZN(_00899_ ) );
INV_X1 _08055_ ( .A(_00715_ ), .ZN(_00900_ ) );
NAND3_X1 _08056_ ( .A1(_00898_ ), .A2(_00899_ ), .A3(_00900_ ), .ZN(_00901_ ) );
OAI21_X1 _08057_ ( .A(\u_idu.imm_branch [2] ), .B1(_00897_ ), .B2(_00901_ ), .ZN(_00902_ ) );
INV_X1 _08058_ ( .A(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00903_ ) );
NAND3_X1 _08059_ ( .A1(_00720_ ), .A2(_00903_ ), .A3(_00677_ ), .ZN(_00904_ ) );
AND2_X2 _08060_ ( .A1(_00902_ ), .A2(_00904_ ), .ZN(_00905_ ) );
INV_X1 _08061_ ( .A(_00905_ ), .ZN(_00906_ ) );
OAI21_X1 _08062_ ( .A(\u_idu.imm_branch [1] ), .B1(_00897_ ), .B2(_00901_ ), .ZN(_00907_ ) );
INV_X1 _08063_ ( .A(_00724_ ), .ZN(_00908_ ) );
OR2_X1 _08064_ ( .A1(_00908_ ), .A2(de_ard_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00909_ ) );
AND2_X2 _08065_ ( .A1(_00907_ ), .A2(_00909_ ), .ZN(_00910_ ) );
INV_X2 _08066_ ( .A(_00910_ ), .ZN(_00911_ ) );
OAI21_X1 _08067_ ( .A(\u_idu.imm_branch [11] ), .B1(_00897_ ), .B2(_00901_ ), .ZN(_00912_ ) );
NAND3_X1 _08068_ ( .A1(_00720_ ), .A2(\u_idu.imm_auipc_lui [12] ), .A3(_00677_ ), .ZN(_00913_ ) );
AND2_X2 _08069_ ( .A1(_00912_ ), .A2(_00913_ ), .ZN(_00914_ ) );
INV_X1 _08070_ ( .A(_00914_ ), .ZN(_00915_ ) );
NAND3_X1 _08071_ ( .A1(_00906_ ), .A2(_00911_ ), .A3(_00915_ ), .ZN(_00916_ ) );
NOR2_X1 _08072_ ( .A1(_00897_ ), .A2(_00901_ ), .ZN(_00917_ ) );
INV_X1 _08073_ ( .A(\u_idu.imm_branch [3] ), .ZN(_00918_ ) );
NOR2_X1 _08074_ ( .A1(_00917_ ), .A2(_00918_ ), .ZN(_00919_ ) );
BUF_X4 _08075_ ( .A(_00919_ ), .Z(_00920_ ) );
AOI21_X4 _08076_ ( .A(_00675_ ), .B1(_00691_ ), .B2(\u_idu.inst [5] ), .ZN(_00921_ ) );
INV_X1 _08077_ ( .A(_00684_ ), .ZN(_00922_ ) );
BUF_X2 _08078_ ( .A(_00922_ ), .Z(_00923_ ) );
AND2_X4 _08079_ ( .A1(_00921_ ), .A2(_00923_ ), .ZN(_00924_ ) );
BUF_X4 _08080_ ( .A(_00924_ ), .Z(_00925_ ) );
NOR2_X2 _08081_ ( .A1(_00925_ ), .A2(_00734_ ), .ZN(_00926_ ) );
NOR2_X2 _08082_ ( .A1(_00924_ ), .A2(_00755_ ), .ZN(_00927_ ) );
BUF_X4 _08083_ ( .A(_00927_ ), .Z(_00928_ ) );
NAND3_X1 _08084_ ( .A1(_00928_ ), .A2(\u_idu.imm_auipc_lui [22] ), .A3(\u_idu.imm_auipc_lui [20] ), .ZN(_00929_ ) );
OAI22_X1 _08085_ ( .A1(_00916_ ), .A2(_00920_ ), .B1(_00926_ ), .B2(_00929_ ), .ZN(_00930_ ) );
NAND4_X1 _08086_ ( .A1(_00898_ ), .A2(_00922_ ), .A3(_00896_ ), .A4(_00899_ ), .ZN(_00931_ ) );
NOR2_X2 _08087_ ( .A1(_00931_ ), .A2(_00691_ ), .ZN(_00932_ ) );
NOR2_X2 _08088_ ( .A1(_00932_ ), .A2(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ), .ZN(_00933_ ) );
AOI21_X1 _08089_ ( .A(_00705_ ), .B1(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ), .B2(_00700_ ), .ZN(_00934_ ) );
NOR2_X4 _08090_ ( .A1(_00933_ ), .A2(_00934_ ), .ZN(_00935_ ) );
OAI21_X1 _08091_ ( .A(\u_idu.imm_auipc_lui [15] ), .B1(_00931_ ), .B2(_00691_ ), .ZN(_00936_ ) );
NAND4_X1 _08092_ ( .A1(_00700_ ), .A2(\u_idu.imm_auipc_lui [15] ), .A3(_00672_ ), .A4(_00703_ ), .ZN(_00937_ ) );
NAND2_X1 _08093_ ( .A1(_00936_ ), .A2(_00937_ ), .ZN(_00938_ ) );
INV_X1 _08094_ ( .A(_00938_ ), .ZN(_00939_ ) );
NOR2_X1 _08095_ ( .A1(_00935_ ), .A2(_00939_ ), .ZN(_00940_ ) );
NAND2_X1 _08096_ ( .A1(_00932_ ), .A2(_00705_ ), .ZN(_00941_ ) );
OAI21_X1 _08097_ ( .A(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_B ), .B1(_00705_ ), .B2(_00700_ ), .ZN(_00942_ ) );
NAND2_X1 _08098_ ( .A1(_00941_ ), .A2(_00942_ ), .ZN(_00943_ ) );
BUF_X4 _08099_ ( .A(_00943_ ), .Z(_00944_ ) );
OAI21_X1 _08100_ ( .A(_00932_ ), .B1(_00718_ ), .B2(_00705_ ), .ZN(_00945_ ) );
INV_X1 _08101_ ( .A(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_1_B ), .ZN(_00946_ ) );
AND2_X1 _08102_ ( .A1(_00945_ ), .A2(_00946_ ), .ZN(_00947_ ) );
BUF_X4 _08103_ ( .A(_00947_ ), .Z(_00948_ ) );
AND3_X1 _08104_ ( .A1(_00940_ ), .A2(_00944_ ), .A3(_00948_ ), .ZN(_00949_ ) );
OAI21_X1 _08105_ ( .A(\u_exu.rlock [7] ), .B1(_00930_ ), .B2(_00949_ ), .ZN(_00950_ ) );
INV_X1 _08106_ ( .A(_00947_ ), .ZN(_00951_ ) );
NAND3_X1 _08107_ ( .A1(_00951_ ), .A2(_00939_ ), .A3(_00935_ ), .ZN(_00952_ ) );
INV_X2 _08108_ ( .A(_00926_ ), .ZN(_00953_ ) );
NOR2_X4 _08109_ ( .A1(_00925_ ), .A2(_00890_ ), .ZN(_00954_ ) );
INV_X1 _08110_ ( .A(_00954_ ), .ZN(_00955_ ) );
INV_X2 _08111_ ( .A(_00927_ ), .ZN(_00956_ ) );
NOR2_X2 _08112_ ( .A1(_00924_ ), .A2(_00748_ ), .ZN(_00957_ ) );
INV_X1 _08113_ ( .A(_00957_ ), .ZN(_00958_ ) );
NAND3_X2 _08114_ ( .A1(_00955_ ), .A2(_00956_ ), .A3(_00958_ ), .ZN(_00959_ ) );
OAI22_X1 _08115_ ( .A1(_00952_ ), .A2(_00943_ ), .B1(_00953_ ), .B2(_00959_ ), .ZN(_00960_ ) );
NAND3_X1 _08116_ ( .A1(_00905_ ), .A2(_00910_ ), .A3(_00914_ ), .ZN(_00961_ ) );
INV_X1 _08117_ ( .A(_00919_ ), .ZN(_00962_ ) );
NOR2_X1 _08118_ ( .A1(_00961_ ), .A2(_00962_ ), .ZN(_00963_ ) );
OAI21_X2 _08119_ ( .A(\u_exu.rlock [8] ), .B1(_00960_ ), .B2(_00963_ ), .ZN(_00964_ ) );
NOR2_X2 _08120_ ( .A1(_00935_ ), .A2(_00938_ ), .ZN(_00965_ ) );
INV_X1 _08121_ ( .A(_00943_ ), .ZN(_00966_ ) );
NAND3_X1 _08122_ ( .A1(_00965_ ), .A2(_00966_ ), .A3(_00947_ ), .ZN(_00967_ ) );
AND2_X4 _08123_ ( .A1(_00928_ ), .A2(_00749_ ), .ZN(_00968_ ) );
NAND3_X1 _08124_ ( .A1(_00968_ ), .A2(\u_idu.imm_auipc_lui [22] ), .A3(_00926_ ), .ZN(_00969_ ) );
NAND2_X1 _08125_ ( .A1(_00967_ ), .A2(_00969_ ), .ZN(_00970_ ) );
NAND3_X1 _08126_ ( .A1(_00906_ ), .A2(_00911_ ), .A3(_00914_ ), .ZN(_00971_ ) );
NOR2_X1 _08127_ ( .A1(_00971_ ), .A2(_00962_ ), .ZN(_00972_ ) );
OAI21_X1 _08128_ ( .A(\u_exu.rlock [14] ), .B1(_00970_ ), .B2(_00972_ ), .ZN(_00973_ ) );
NAND2_X1 _08129_ ( .A1(_00964_ ), .A2(_00973_ ), .ZN(_00974_ ) );
AND2_X2 _08130_ ( .A1(_00935_ ), .A2(_00938_ ), .ZN(_00975_ ) );
BUF_X4 _08131_ ( .A(_00975_ ), .Z(_00976_ ) );
NAND3_X1 _08132_ ( .A1(_00976_ ), .A2(_00943_ ), .A3(_00948_ ), .ZN(_00977_ ) );
BUF_X2 _08133_ ( .A(_00755_ ), .Z(_00978_ ) );
AND2_X1 _08134_ ( .A1(_00957_ ), .A2(_00978_ ), .ZN(_00979_ ) );
BUF_X4 _08135_ ( .A(_00979_ ), .Z(_00980_ ) );
NAND3_X1 _08136_ ( .A1(_00980_ ), .A2(\u_idu.imm_auipc_lui [22] ), .A3(_00953_ ), .ZN(_00981_ ) );
NAND3_X1 _08137_ ( .A1(_00906_ ), .A2(_00915_ ), .A3(_00910_ ), .ZN(_00982_ ) );
OAI211_X1 _08138_ ( .A(_00977_ ), .B(_00981_ ), .C1(_00919_ ), .C2(_00982_ ), .ZN(_00983_ ) );
OAI22_X1 _08139_ ( .A1(_00952_ ), .A2(_00966_ ), .B1(_00926_ ), .B2(_00959_ ), .ZN(_00984_ ) );
NOR2_X1 _08140_ ( .A1(_00961_ ), .A2(_00919_ ), .ZN(_00985_ ) );
OR2_X1 _08141_ ( .A1(_00984_ ), .A2(_00985_ ), .ZN(_00986_ ) );
AOI221_X2 _08142_ ( .A(_00974_ ), .B1(\u_exu.rlock [5] ), .B2(_00983_ ), .C1(\u_exu.rlock [0] ), .C2(_00986_ ), .ZN(_00987_ ) );
NAND3_X1 _08143_ ( .A1(_00976_ ), .A2(_00966_ ), .A3(_00951_ ), .ZN(_00988_ ) );
BUF_X2 _08144_ ( .A(_00957_ ), .Z(_00989_ ) );
NAND3_X1 _08145_ ( .A1(_00989_ ), .A2(_00890_ ), .A3(_00978_ ), .ZN(_00990_ ) );
OAI21_X1 _08146_ ( .A(_00988_ ), .B1(_00888_ ), .B2(_00990_ ), .ZN(_00991_ ) );
NAND3_X1 _08147_ ( .A1(_00915_ ), .A2(_00905_ ), .A3(_00910_ ), .ZN(_00992_ ) );
BUF_X4 _08148_ ( .A(_00962_ ), .Z(_00993_ ) );
NOR2_X1 _08149_ ( .A1(_00992_ ), .A2(_00993_ ), .ZN(_00994_ ) );
OAI21_X1 _08150_ ( .A(\u_exu.rlock [9] ), .B1(_00991_ ), .B2(_00994_ ), .ZN(_00995_ ) );
NAND3_X1 _08151_ ( .A1(_00976_ ), .A2(_00966_ ), .A3(_00948_ ), .ZN(_00996_ ) );
NAND3_X1 _08152_ ( .A1(_00980_ ), .A2(\u_idu.imm_auipc_lui [22] ), .A3(_00926_ ), .ZN(_00997_ ) );
NAND2_X1 _08153_ ( .A1(_00996_ ), .A2(_00997_ ), .ZN(_00998_ ) );
NOR2_X1 _08154_ ( .A1(_00982_ ), .A2(_00993_ ), .ZN(_00999_ ) );
OAI21_X1 _08155_ ( .A(\u_exu.rlock [13] ), .B1(_00998_ ), .B2(_00999_ ), .ZN(_01000_ ) );
AND2_X1 _08156_ ( .A1(_00995_ ), .A2(_01000_ ), .ZN(_01001_ ) );
OAI22_X1 _08157_ ( .A1(_00916_ ), .A2(_00993_ ), .B1(_00953_ ), .B2(_00929_ ), .ZN(_01002_ ) );
AND3_X1 _08158_ ( .A1(_00940_ ), .A2(_00966_ ), .A3(_00948_ ), .ZN(_01003_ ) );
OAI21_X1 _08159_ ( .A(\u_exu.rlock [15] ), .B1(_01002_ ), .B2(_01003_ ), .ZN(_01004_ ) );
NAND3_X1 _08160_ ( .A1(_00940_ ), .A2(_00951_ ), .A3(_00944_ ), .ZN(_01005_ ) );
NAND4_X1 _08161_ ( .A1(_00957_ ), .A2(_00888_ ), .A3(_00890_ ), .A4(fanout_net_20 ), .ZN(_01006_ ) );
NAND2_X1 _08162_ ( .A1(_01005_ ), .A2(_01006_ ), .ZN(_01007_ ) );
NAND3_X1 _08163_ ( .A1(_00911_ ), .A2(_00915_ ), .A3(_00905_ ), .ZN(_01008_ ) );
NOR2_X1 _08164_ ( .A1(_01008_ ), .A2(_00920_ ), .ZN(_01009_ ) );
OAI21_X1 _08165_ ( .A(\u_exu.rlock [3] ), .B1(_01007_ ), .B2(_01009_ ), .ZN(_01010_ ) );
AND3_X1 _08166_ ( .A1(_00965_ ), .A2(_00951_ ), .A3(_00966_ ), .ZN(_01011_ ) );
NAND3_X1 _08167_ ( .A1(_00968_ ), .A2(_00890_ ), .A3(_00926_ ), .ZN(_01012_ ) );
NAND3_X1 _08168_ ( .A1(_00911_ ), .A2(_00905_ ), .A3(_00914_ ), .ZN(_01013_ ) );
OAI21_X1 _08169_ ( .A(_01012_ ), .B1(_01013_ ), .B2(_00993_ ), .ZN(_01014_ ) );
OAI21_X1 _08170_ ( .A(\u_exu.rlock [10] ), .B1(_01011_ ), .B2(_01014_ ), .ZN(_01015_ ) );
AND2_X2 _08171_ ( .A1(_00935_ ), .A2(_00939_ ), .ZN(_01016_ ) );
BUF_X4 _08172_ ( .A(_01016_ ), .Z(_01017_ ) );
AND3_X1 _08173_ ( .A1(_01017_ ), .A2(_00966_ ), .A3(_00948_ ), .ZN(_01018_ ) );
NOR2_X1 _08174_ ( .A1(_00928_ ), .A2(_00957_ ), .ZN(_01019_ ) );
NAND3_X1 _08175_ ( .A1(_01019_ ), .A2(_00954_ ), .A3(_00926_ ), .ZN(_01020_ ) );
NAND3_X1 _08176_ ( .A1(_00906_ ), .A2(_00910_ ), .A3(_00914_ ), .ZN(_01021_ ) );
OAI21_X1 _08177_ ( .A(_01020_ ), .B1(_01021_ ), .B2(_00993_ ), .ZN(_01022_ ) );
OAI21_X1 _08178_ ( .A(\u_exu.rlock [12] ), .B1(_01018_ ), .B2(_01022_ ), .ZN(_01023_ ) );
AND4_X1 _08179_ ( .A1(_01004_ ), .A2(_01010_ ), .A3(_01015_ ), .A4(_01023_ ), .ZN(_01024_ ) );
AND4_X2 _08180_ ( .A1(_00950_ ), .A2(_00987_ ), .A3(_01001_ ), .A4(_01024_ ), .ZN(_01025_ ) );
BUF_X4 _08181_ ( .A(_00951_ ), .Z(_01026_ ) );
NAND3_X1 _08182_ ( .A1(_00965_ ), .A2(_01026_ ), .A3(_00944_ ), .ZN(_01027_ ) );
BUF_X2 _08183_ ( .A(_00953_ ), .Z(_01028_ ) );
NAND3_X1 _08184_ ( .A1(_00968_ ), .A2(_00890_ ), .A3(_01028_ ), .ZN(_01029_ ) );
NAND2_X1 _08185_ ( .A1(_01027_ ), .A2(_01029_ ), .ZN(_01030_ ) );
NOR2_X1 _08186_ ( .A1(_01013_ ), .A2(_00920_ ), .ZN(_01031_ ) );
OAI21_X1 _08187_ ( .A(\u_exu.rlock [2] ), .B1(_01030_ ), .B2(_01031_ ), .ZN(_01032_ ) );
NAND3_X1 _08188_ ( .A1(_00965_ ), .A2(_00944_ ), .A3(_00948_ ), .ZN(_01033_ ) );
NAND3_X1 _08189_ ( .A1(_00968_ ), .A2(\u_idu.imm_auipc_lui [22] ), .A3(_00953_ ), .ZN(_01034_ ) );
NAND2_X1 _08190_ ( .A1(_01033_ ), .A2(_01034_ ), .ZN(_01035_ ) );
NOR2_X1 _08191_ ( .A1(_00971_ ), .A2(_00920_ ), .ZN(_01036_ ) );
OAI21_X1 _08192_ ( .A(\u_exu.rlock [6] ), .B1(_01035_ ), .B2(_01036_ ), .ZN(_01037_ ) );
AND3_X1 _08193_ ( .A1(_00976_ ), .A2(_00944_ ), .A3(_01026_ ), .ZN(_01038_ ) );
OAI22_X1 _08194_ ( .A1(_00992_ ), .A2(_00920_ ), .B1(\u_idu.imm_auipc_lui [23] ), .B2(_00990_ ), .ZN(_01039_ ) );
OAI21_X2 _08195_ ( .A(\u_exu.rlock [1] ), .B1(_01038_ ), .B2(_01039_ ), .ZN(_01040_ ) );
NAND4_X1 _08196_ ( .A1(_00989_ ), .A2(\u_idu.imm_auipc_lui [23] ), .A3(_00890_ ), .A4(fanout_net_20 ), .ZN(_01041_ ) );
OAI21_X1 _08197_ ( .A(_01041_ ), .B1(_01008_ ), .B2(_00993_ ), .ZN(_01042_ ) );
BUF_X2 _08198_ ( .A(_00966_ ), .Z(_01043_ ) );
AND3_X1 _08199_ ( .A1(_00940_ ), .A2(_01026_ ), .A3(_01043_ ), .ZN(_01044_ ) );
OAI21_X1 _08200_ ( .A(\u_exu.rlock [11] ), .B1(_01042_ ), .B2(_01044_ ), .ZN(_01045_ ) );
NAND4_X1 _08201_ ( .A1(_01032_ ), .A2(_01037_ ), .A3(_01040_ ), .A4(_01045_ ), .ZN(_01046_ ) );
INV_X1 _08202_ ( .A(\u_exu.rlock [4] ), .ZN(_01047_ ) );
NOR2_X1 _08203_ ( .A1(_01021_ ), .A2(_00920_ ), .ZN(_01048_ ) );
BUF_X4 _08204_ ( .A(_00954_ ), .Z(_01049_ ) );
AND3_X1 _08205_ ( .A1(_01019_ ), .A2(_01049_ ), .A3(_00953_ ), .ZN(_01050_ ) );
NOR2_X1 _08206_ ( .A1(_01048_ ), .A2(_01050_ ), .ZN(_01051_ ) );
NAND3_X1 _08207_ ( .A1(_01017_ ), .A2(_00944_ ), .A3(_00948_ ), .ZN(_01052_ ) );
AOI21_X1 _08208_ ( .A(_01047_ ), .B1(_01051_ ), .B2(_01052_ ), .ZN(_01053_ ) );
NOR4_X2 _08209_ ( .A1(_01046_ ), .A2(\u_exu.exe_start ), .A3(_00767_ ), .A4(_01053_ ), .ZN(_01054_ ) );
AND2_X2 _08210_ ( .A1(_01025_ ), .A2(_01054_ ), .ZN(_01055_ ) );
INV_X4 _08211_ ( .A(_01055_ ), .ZN(_01056_ ) );
BUF_X4 _08212_ ( .A(_01056_ ), .Z(_01057_ ) );
NOR2_X1 _08213_ ( .A1(_00695_ ), .A2(\u_idu.imm_auipc_lui [14] ), .ZN(_01058_ ) );
NOR2_X1 _08214_ ( .A1(\u_idu.imm_auipc_lui [13] ), .A2(\u_exu.alu_ctrl_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A ), .ZN(_01059_ ) );
OAI21_X1 _08215_ ( .A(_00711_ ), .B1(_01058_ ), .B2(_01059_ ), .ZN(_01060_ ) );
AOI21_X1 _08216_ ( .A(_00896_ ), .B1(_00668_ ), .B2(_00652_ ), .ZN(_01061_ ) );
NOR2_X1 _08217_ ( .A1(_01061_ ), .A2(_00687_ ), .ZN(_01062_ ) );
AOI211_X1 _08218_ ( .A(_00894_ ), .B(_01057_ ), .C1(_01060_ ), .C2(_01062_ ), .ZN(_00122_ ) );
NOR3_X1 _08219_ ( .A1(_01058_ ), .A2(_00903_ ), .A3(\u_idu.imm_auipc_lui [12] ), .ZN(_01063_ ) );
AOI21_X1 _08220_ ( .A(\u_idu.imm_auipc_lui [13] ), .B1(_00646_ ), .B2(\u_idu.imm_auipc_lui [14] ), .ZN(_01064_ ) );
OR3_X1 _08221_ ( .A1(_00898_ ), .A2(_01063_ ), .A3(_01064_ ), .ZN(_01065_ ) );
NOR2_X1 _08222_ ( .A1(_00660_ ), .A2(_00896_ ), .ZN(_01066_ ) );
AND2_X1 _08223_ ( .A1(_00704_ ), .A2(_00697_ ), .ZN(_01067_ ) );
NOR3_X1 _08224_ ( .A1(_01066_ ), .A2(_00687_ ), .A3(_01067_ ), .ZN(_01068_ ) );
AOI211_X1 _08225_ ( .A(_00894_ ), .B(_01057_ ), .C1(_01065_ ), .C2(_01068_ ), .ZN(_00123_ ) );
NOR2_X1 _08226_ ( .A1(_01055_ ), .A2(_00892_ ), .ZN(_01069_ ) );
BUF_X2 _08227_ ( .A(_01069_ ), .Z(_01070_ ) );
NOR2_X1 _08228_ ( .A1(_00744_ ), .A2(_00680_ ), .ZN(_01071_ ) );
AND4_X1 _08229_ ( .A1(_00648_ ), .A2(_00672_ ), .A3(_00665_ ), .A4(_00703_ ), .ZN(_01072_ ) );
AOI21_X1 _08230_ ( .A(_01072_ ), .B1(_00692_ ), .B2(_00701_ ), .ZN(_01073_ ) );
NAND2_X1 _08231_ ( .A1(_01071_ ), .A2(_01073_ ), .ZN(_01074_ ) );
AND2_X1 _08232_ ( .A1(_00713_ ), .A2(_00710_ ), .ZN(_01075_ ) );
NOR2_X1 _08233_ ( .A1(_01074_ ), .A2(_01075_ ), .ZN(_01076_ ) );
AND2_X1 _08234_ ( .A1(\u_idu.inst [5] ), .A2(\u_idu.inst [4] ), .ZN(_01077_ ) );
AND2_X1 _08235_ ( .A1(_00689_ ), .A2(_01077_ ), .ZN(_01078_ ) );
NAND2_X1 _08236_ ( .A1(_00664_ ), .A2(_00658_ ), .ZN(_01079_ ) );
AND2_X1 _08237_ ( .A1(_00667_ ), .A2(_00860_ ), .ZN(_01080_ ) );
OAI21_X1 _08238_ ( .A(_01078_ ), .B1(_01079_ ), .B2(_01080_ ), .ZN(_01081_ ) );
AND2_X1 _08239_ ( .A1(_00655_ ), .A2(\u_idu.imm_auipc_lui [14] ), .ZN(_01082_ ) );
NAND2_X1 _08240_ ( .A1(\u_idu.imm_auipc_lui [12] ), .A2(\u_idu.imm_auipc_lui [14] ), .ZN(_01083_ ) );
NOR2_X1 _08241_ ( .A1(_01083_ ), .A2(\u_idu.imm_auipc_lui [13] ), .ZN(_01084_ ) );
OR2_X1 _08242_ ( .A1(_01082_ ), .A2(_01084_ ), .ZN(_01085_ ) );
OAI21_X1 _08243_ ( .A(_00711_ ), .B1(_01085_ ), .B2(_01063_ ), .ZN(_01086_ ) );
OAI21_X1 _08244_ ( .A(_00684_ ), .B1(_00693_ ), .B2(_00718_ ), .ZN(_01087_ ) );
AND3_X1 _08245_ ( .A1(_01081_ ), .A2(_01086_ ), .A3(_01087_ ), .ZN(_01088_ ) );
AOI211_X1 _08246_ ( .A(_00764_ ), .B(_00879_ ), .C1(_01076_ ), .C2(_01088_ ), .ZN(_01089_ ) );
OR2_X1 _08247_ ( .A1(_01070_ ), .A2(_01089_ ), .ZN(_00124_ ) );
BUF_X2 _08248_ ( .A(_01055_ ), .Z(_01090_ ) );
AOI211_X1 _08249_ ( .A(_00764_ ), .B(_00879_ ), .C1(_01071_ ), .C2(_00758_ ), .ZN(_00231_ ) );
INV_X1 _08250_ ( .A(_00691_ ), .ZN(_01091_ ) );
NOR3_X1 _08251_ ( .A1(_01091_ ), .A2(_00682_ ), .A3(_00706_ ), .ZN(_01092_ ) );
INV_X1 _08252_ ( .A(_00678_ ), .ZN(_01093_ ) );
NOR2_X1 _08253_ ( .A1(_00693_ ), .A2(_01084_ ), .ZN(_01094_ ) );
AOI21_X1 _08254_ ( .A(_01093_ ), .B1(_01094_ ), .B2(_00698_ ), .ZN(_01095_ ) );
NOR3_X1 _08255_ ( .A1(_01092_ ), .A2(_01095_ ), .A3(_00707_ ), .ZN(_01096_ ) );
AND4_X1 _08256_ ( .A1(_00749_ ), .A2(_00754_ ), .A3(_00732_ ), .A4(_00731_ ), .ZN(_01097_ ) );
AND4_X1 _08257_ ( .A1(_00888_ ), .A2(_01097_ ), .A3(_00704_ ), .A4(_00756_ ), .ZN(_01098_ ) );
NAND2_X1 _08258_ ( .A1(_01098_ ), .A2(_00718_ ), .ZN(_01099_ ) );
AND2_X1 _08259_ ( .A1(_01096_ ), .A2(_01099_ ), .ZN(_01100_ ) );
AND3_X1 _08260_ ( .A1(_00692_ ), .A2(_00646_ ), .A3(_00648_ ), .ZN(_01101_ ) );
OAI211_X1 _08261_ ( .A(_00646_ ), .B(_00695_ ), .C1(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .C2(\u_idu.imm_auipc_lui [14] ), .ZN(_01102_ ) );
AOI21_X1 _08262_ ( .A(_01093_ ), .B1(_00698_ ), .B2(_01102_ ), .ZN(_01103_ ) );
NOR3_X1 _08263_ ( .A1(_01101_ ), .A2(_00707_ ), .A3(_01103_ ), .ZN(_01104_ ) );
AND4_X1 _08264_ ( .A1(_01090_ ), .A2(_00231_ ), .A3(_01100_ ), .A4(_01104_ ), .ZN(_00125_ ) );
BUF_X4 _08265_ ( .A(_01025_ ), .Z(_01105_ ) );
BUF_X8 _08266_ ( .A(_01105_ ), .Z(_01106_ ) );
BUF_X8 _08267_ ( .A(_01106_ ), .Z(_01107_ ) );
BUF_X4 _08268_ ( .A(_01054_ ), .Z(_01108_ ) );
BUF_X4 _08269_ ( .A(_01108_ ), .Z(_01109_ ) );
CLKBUF_X2 _08270_ ( .A(_01109_ ), .Z(_01110_ ) );
AOI21_X1 _08271_ ( .A(_00688_ ), .B1(_00694_ ), .B2(_01083_ ), .ZN(_01111_ ) );
NOR2_X1 _08272_ ( .A1(_01111_ ), .A2(_00725_ ), .ZN(_01112_ ) );
NAND3_X1 _08273_ ( .A1(_01097_ ), .A2(_00888_ ), .A3(_00756_ ), .ZN(_01113_ ) );
NAND4_X1 _08274_ ( .A1(_00730_ ), .A2(_00733_ ), .A3(_00888_ ), .A4(_00749_ ), .ZN(_01114_ ) );
AOI21_X1 _08275_ ( .A(_00700_ ), .B1(_01113_ ), .B2(_01114_ ), .ZN(_01115_ ) );
NAND2_X1 _08276_ ( .A1(_00875_ ), .A2(_00706_ ), .ZN(_01116_ ) );
OAI21_X1 _08277_ ( .A(_00704_ ), .B1(_01115_ ), .B2(_01116_ ), .ZN(_01117_ ) );
AND2_X1 _08278_ ( .A1(_01112_ ), .A2(_01117_ ), .ZN(_01118_ ) );
NOR3_X1 _08279_ ( .A1(_01118_ ), .A2(_00855_ ), .A3(_00879_ ), .ZN(_00229_ ) );
AND3_X1 _08280_ ( .A1(_01107_ ), .A2(_01110_ ), .A3(_00229_ ), .ZN(_00126_ ) );
AND3_X1 _08281_ ( .A1(_00667_ ), .A2(_00860_ ), .A3(\u_idu.imm_auipc_lui [30] ), .ZN(_01119_ ) );
AND2_X1 _08282_ ( .A1(_00647_ ), .A2(_00651_ ), .ZN(_01120_ ) );
OAI21_X1 _08283_ ( .A(_00675_ ), .B1(_01119_ ), .B2(_01120_ ), .ZN(_01121_ ) );
OAI21_X1 _08284_ ( .A(_00678_ ), .B1(_00693_ ), .B2(_00718_ ), .ZN(_01122_ ) );
NAND2_X1 _08285_ ( .A1(_00684_ ), .A2(_01085_ ), .ZN(_01123_ ) );
NAND4_X1 _08286_ ( .A1(_00672_ ), .A2(_00646_ ), .A3(_00710_ ), .A4(_01058_ ), .ZN(_01124_ ) );
NAND4_X1 _08287_ ( .A1(_01121_ ), .A2(_01122_ ), .A3(_01123_ ), .A4(_01124_ ), .ZN(_01125_ ) );
NOR4_X1 _08288_ ( .A1(_00898_ ), .A2(\u_idu.imm_auipc_lui [13] ), .A3(\u_exu.opt_$_NOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B ), .A4(_01083_ ), .ZN(_01126_ ) );
OAI211_X1 _08289_ ( .A(_00865_ ), .B(_00862_ ), .C1(_01125_ ), .C2(_01126_ ), .ZN(_01127_ ) );
INV_X1 _08290_ ( .A(_01127_ ), .ZN(_00230_ ) );
AND3_X1 _08291_ ( .A1(_01107_ ), .A2(_01110_ ), .A3(_00230_ ), .ZN(_00127_ ) );
NOR3_X1 _08292_ ( .A1(_00695_ ), .A2(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(\u_idu.imm_auipc_lui [12] ), .ZN(_01128_ ) );
OAI21_X1 _08293_ ( .A(_00711_ ), .B1(_01058_ ), .B2(_01128_ ), .ZN(_01129_ ) );
NAND3_X1 _08294_ ( .A1(_00661_ ), .A2(_00860_ ), .A3(\u_idu.imm_auipc_lui [30] ), .ZN(_01130_ ) );
AOI21_X1 _08295_ ( .A(_00896_ ), .B1(_00653_ ), .B2(_01130_ ), .ZN(_01131_ ) );
NOR3_X1 _08296_ ( .A1(_01131_ ), .A2(_00687_ ), .A3(_01067_ ), .ZN(_01132_ ) );
AOI211_X1 _08297_ ( .A(_00894_ ), .B(_01057_ ), .C1(_01129_ ), .C2(_01132_ ), .ZN(_00128_ ) );
AND3_X1 _08298_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [31] ), .ZN(_01133_ ) );
NAND2_X1 _08299_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .ZN(_01134_ ) );
BUF_X4 _08300_ ( .A(_01134_ ), .Z(_01135_ ) );
BUF_X4 _08301_ ( .A(_01135_ ), .Z(_01136_ ) );
AOI211_X1 _08302_ ( .A(fanout_net_9 ), .B(_01133_ ), .C1(\ea_addr [31] ), .C2(_01136_ ), .ZN(_01137_ ) );
INV_X32 _08303_ ( .A(icah_valid ), .ZN(_01138_ ) );
NOR2_X4 _08304_ ( .A1(_01138_ ), .A2(\u_arbiter.working ), .ZN(_01139_ ) );
BUF_X8 _08305_ ( .A(_01139_ ), .Z(_01140_ ) );
INV_X1 _08306_ ( .A(\u_arbiter.raddr [0] ), .ZN(_01141_ ) );
NOR2_X2 _08307_ ( .A1(_01140_ ), .A2(_01141_ ), .ZN(\io_master_araddr [0] ) );
INV_X1 _08308_ ( .A(\u_arbiter.raddr [1] ), .ZN(_01142_ ) );
AND2_X2 _08309_ ( .A1(\io_master_araddr [0] ), .A2(_01142_ ), .ZN(_01143_ ) );
INV_X2 _08310_ ( .A(_01143_ ), .ZN(_01144_ ) );
BUF_X8 _08311_ ( .A(_01139_ ), .Z(_01145_ ) );
MUX2_X1 _08312_ ( .A(\u_arbiter.raddr [22] ), .B(\ca_addr [22] ), .S(_01145_ ), .Z(\io_master_araddr [22] ) );
MUX2_X1 _08313_ ( .A(\u_arbiter.raddr [17] ), .B(\ca_addr [17] ), .S(_01140_ ), .Z(\io_master_araddr [17] ) );
NOR2_X1 _08314_ ( .A1(\io_master_araddr [22] ), .A2(\io_master_araddr [17] ), .ZN(_01146_ ) );
MUX2_X1 _08315_ ( .A(\u_arbiter.raddr [21] ), .B(\ca_addr [21] ), .S(_01140_ ), .Z(\io_master_araddr [21] ) );
BUF_X32 _08316_ ( .A(_00634_ ), .Z(_01147_ ) );
AND3_X1 _08317_ ( .A1(_01147_ ), .A2(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_B ), .A3(icah_valid ), .ZN(_01148_ ) );
INV_X1 _08318_ ( .A(_01145_ ), .ZN(_01149_ ) );
AOI21_X4 _08319_ ( .A(_01148_ ), .B1(_01149_ ), .B2(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_A ), .ZN(\io_master_araddr [18] ) );
NOR2_X1 _08320_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [18] ), .ZN(_01150_ ) );
NAND2_X1 _08321_ ( .A1(_01146_ ), .A2(_01150_ ), .ZN(_01151_ ) );
MUX2_X1 _08322_ ( .A(\u_arbiter.raddr [19] ), .B(\ca_addr [19] ), .S(_01140_ ), .Z(\io_master_araddr [19] ) );
OAI21_X1 _08323_ ( .A(\u_arbiter.raddr [16] ), .B1(_01138_ ), .B2(\u_arbiter.working ), .ZN(_01152_ ) );
OAI21_X1 _08324_ ( .A(\u_arbiter.raddr [23] ), .B1(_01138_ ), .B2(\u_arbiter.working ), .ZN(_01153_ ) );
NAND3_X1 _08325_ ( .A1(_01147_ ), .A2(\ca_addr [16] ), .A3(icah_valid ), .ZN(_01154_ ) );
NAND3_X1 _08326_ ( .A1(_01147_ ), .A2(\ca_addr [23] ), .A3(icah_valid ), .ZN(_01155_ ) );
NAND4_X2 _08327_ ( .A1(_01152_ ), .A2(_01153_ ), .A3(_01154_ ), .A4(_01155_ ), .ZN(_01156_ ) );
OAI21_X1 _08328_ ( .A(\u_arbiter.raddr [20] ), .B1(_01138_ ), .B2(\u_arbiter.working ), .ZN(_01157_ ) );
NAND3_X1 _08329_ ( .A1(_01147_ ), .A2(\ca_addr [20] ), .A3(icah_valid ), .ZN(_01158_ ) );
NAND2_X1 _08330_ ( .A1(_01157_ ), .A2(_01158_ ), .ZN(\io_master_araddr [20] ) );
OR3_X4 _08331_ ( .A1(\io_master_araddr [19] ), .A2(_01156_ ), .A3(\io_master_araddr [20] ), .ZN(_01159_ ) );
NOR2_X2 _08332_ ( .A1(_01151_ ), .A2(_01159_ ), .ZN(_01160_ ) );
NOR3_X1 _08333_ ( .A1(_01138_ ), .A2(\ca_addr [9] ), .A3(\u_arbiter.working ), .ZN(_01161_ ) );
AOI21_X2 _08334_ ( .A(\u_arbiter.raddr [9] ), .B1(_01147_ ), .B2(icah_valid ), .ZN(_01162_ ) );
NOR2_X1 _08335_ ( .A1(_01161_ ), .A2(_01162_ ), .ZN(\io_master_araddr [9] ) );
OAI21_X1 _08336_ ( .A(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_A ), .B1(_01138_ ), .B2(\u_arbiter.working ), .ZN(_01163_ ) );
NAND3_X2 _08337_ ( .A1(_01147_ ), .A2(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_B ), .A3(icah_valid ), .ZN(_01164_ ) );
AND2_X2 _08338_ ( .A1(_01163_ ), .A2(_01164_ ), .ZN(\io_master_araddr [10] ) );
OAI21_X1 _08339_ ( .A(\u_arbiter.raddr [13] ), .B1(_01138_ ), .B2(\u_arbiter.working ), .ZN(_01165_ ) );
NAND3_X1 _08340_ ( .A1(_01147_ ), .A2(\ca_addr [13] ), .A3(icah_valid ), .ZN(_01166_ ) );
NAND2_X1 _08341_ ( .A1(_01165_ ), .A2(_01166_ ), .ZN(\io_master_araddr [13] ) );
OAI21_X2 _08342_ ( .A(\u_arbiter.raddr [12] ), .B1(_01138_ ), .B2(\u_arbiter.working ), .ZN(_01167_ ) );
NAND3_X2 _08343_ ( .A1(_01147_ ), .A2(\ca_addr [12] ), .A3(icah_valid ), .ZN(_01168_ ) );
NAND2_X2 _08344_ ( .A1(_01167_ ), .A2(_01168_ ), .ZN(\io_master_araddr [12] ) );
OR4_X4 _08345_ ( .A1(\io_master_araddr [9] ), .A2(\io_master_araddr [10] ), .A3(\io_master_araddr [13] ), .A4(\io_master_araddr [12] ), .ZN(_01169_ ) );
BUF_X32 _08346_ ( .A(_01138_ ), .Z(_01170_ ) );
OR3_X4 _08347_ ( .A1(_01170_ ), .A2(\u_arbiter.working ), .A3(\u_icache.caddr_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ), .ZN(_01171_ ) );
AOI21_X1 _08348_ ( .A(\u_arbiter.raddr [14] ), .B1(_00635_ ), .B2(icah_valid ), .ZN(_01172_ ) );
NOR3_X1 _08349_ ( .A1(_01170_ ), .A2(\ca_addr [14] ), .A3(\u_arbiter.working ), .ZN(_01173_ ) );
OAI221_X1 _08350_ ( .A(_01171_ ), .B1(\u_icache.caddr_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_MUX__B_A ), .B2(_01145_ ), .C1(_01172_ ), .C2(_01173_ ), .ZN(_01174_ ) );
NOR2_X4 _08351_ ( .A1(_01169_ ), .A2(_01174_ ), .ZN(_01175_ ) );
MUX2_X1 _08352_ ( .A(\u_arbiter.raddr [24] ), .B(\ca_addr [24] ), .S(_01140_ ), .Z(\io_master_araddr [24] ) );
MUX2_X1 _08353_ ( .A(\u_arbiter.raddr [25] ), .B(\ca_addr [25] ), .S(_01140_ ), .Z(\io_master_araddr [25] ) );
NOR2_X1 _08354_ ( .A1(\io_master_araddr [24] ), .A2(\io_master_araddr [25] ), .ZN(_01176_ ) );
MUX2_X1 _08355_ ( .A(\u_arbiter.raddr [11] ), .B(\ca_addr [11] ), .S(_01140_ ), .Z(\io_master_araddr [11] ) );
MUX2_X1 _08356_ ( .A(\u_arbiter.raddr [15] ), .B(\ca_addr [15] ), .S(_01140_ ), .Z(\io_master_araddr [15] ) );
NOR2_X1 _08357_ ( .A1(\io_master_araddr [11] ), .A2(\io_master_araddr [15] ), .ZN(_01177_ ) );
MUX2_X1 _08358_ ( .A(\u_arbiter.raddr [27] ), .B(\ca_addr [27] ), .S(_01140_ ), .Z(\io_master_araddr [27] ) );
INV_X1 _08359_ ( .A(io_master_araddr_$_NOT__Y_5_A_$_MUX__Y_B ), .ZN(_01178_ ) );
NAND3_X1 _08360_ ( .A1(_01178_ ), .A2(_01147_ ), .A3(icah_valid ), .ZN(_01179_ ) );
OAI21_X1 _08361_ ( .A(_01179_ ), .B1(_01145_ ), .B2(io_master_araddr_$_NOT__Y_5_A_$_MUX__Y_A ), .ZN(\io_master_araddr [26] ) );
NOR2_X1 _08362_ ( .A1(\io_master_araddr [27] ), .A2(\io_master_araddr [26] ), .ZN(_01180_ ) );
AND3_X1 _08363_ ( .A1(_01176_ ), .A2(_01177_ ), .A3(_01180_ ), .ZN(_01181_ ) );
AND3_X1 _08364_ ( .A1(_01160_ ), .A2(_01175_ ), .A3(_01181_ ), .ZN(_01182_ ) );
OAI21_X2 _08365_ ( .A(\u_arbiter.raddr [7] ), .B1(_01170_ ), .B2(\u_arbiter.working ), .ZN(_01183_ ) );
NAND3_X1 _08366_ ( .A1(_00635_ ), .A2(\ca_addr [7] ), .A3(icah_valid ), .ZN(_01184_ ) );
NAND2_X1 _08367_ ( .A1(_01183_ ), .A2(_01184_ ), .ZN(\io_master_araddr [7] ) );
INV_X1 _08368_ ( .A(\io_master_araddr [7] ), .ZN(_01185_ ) );
MUX2_X1 _08369_ ( .A(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_A ), .B(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_B ), .S(_01145_ ), .Z(_01186_ ) );
INV_X1 _08370_ ( .A(_01186_ ), .ZN(\io_master_araddr [4] ) );
MUX2_X1 _08371_ ( .A(\u_arbiter.raddr [5] ), .B(\ca_addr [5] ), .S(_01145_ ), .Z(\io_master_araddr [5] ) );
NOR2_X1 _08372_ ( .A1(\io_master_araddr [4] ), .A2(\io_master_araddr [5] ), .ZN(_01187_ ) );
OAI21_X2 _08373_ ( .A(\u_icache.caddr_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_MUX__B_A ), .B1(_01170_ ), .B2(\u_arbiter.working ), .ZN(_01188_ ) );
NAND3_X1 _08374_ ( .A1(_00635_ ), .A2(icah_valid ), .A3(\u_icache.caddr_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ), .ZN(_01189_ ) );
AND2_X2 _08375_ ( .A1(_01188_ ), .A2(_01189_ ), .ZN(\io_master_araddr [6] ) );
NAND2_X1 _08376_ ( .A1(_01185_ ), .A2(\io_master_araddr [6] ), .ZN(_01190_ ) );
OAI211_X1 _08377_ ( .A(_01182_ ), .B(_01185_ ), .C1(_01187_ ), .C2(_01190_ ), .ZN(_01191_ ) );
NOR3_X1 _08378_ ( .A1(_01170_ ), .A2(\ca_addr [28] ), .A3(\u_arbiter.working ), .ZN(_01192_ ) );
AOI21_X2 _08379_ ( .A(\u_arbiter.raddr [28] ), .B1(_00635_ ), .B2(icah_valid ), .ZN(_01193_ ) );
NOR2_X1 _08380_ ( .A1(_01192_ ), .A2(_01193_ ), .ZN(\io_master_araddr [28] ) );
OAI21_X2 _08381_ ( .A(\u_arbiter.raddr [30] ), .B1(_01170_ ), .B2(\u_arbiter.working ), .ZN(_01194_ ) );
NAND3_X1 _08382_ ( .A1(_00635_ ), .A2(\ca_addr [30] ), .A3(icah_valid ), .ZN(_01195_ ) );
NAND2_X1 _08383_ ( .A1(_01194_ ), .A2(_01195_ ), .ZN(\io_master_araddr [30] ) );
NOR2_X1 _08384_ ( .A1(\io_master_araddr [28] ), .A2(\io_master_araddr [30] ), .ZN(_01196_ ) );
OAI21_X1 _08385_ ( .A(\u_arbiter.raddr [31] ), .B1(_01170_ ), .B2(\u_arbiter.working ), .ZN(_01197_ ) );
NAND3_X1 _08386_ ( .A1(_00635_ ), .A2(\ca_addr [31] ), .A3(icah_valid ), .ZN(_01198_ ) );
OAI21_X1 _08387_ ( .A(\u_arbiter.raddr [29] ), .B1(_01170_ ), .B2(\u_arbiter.working ), .ZN(_01199_ ) );
NAND3_X1 _08388_ ( .A1(_00635_ ), .A2(\ca_addr [29] ), .A3(icah_valid ), .ZN(_01200_ ) );
AOI22_X1 _08389_ ( .A1(_01197_ ), .A2(_01198_ ), .B1(_01199_ ), .B2(_01200_ ), .ZN(_01201_ ) );
AND2_X4 _08390_ ( .A1(_01196_ ), .A2(_01201_ ), .ZN(_01202_ ) );
NAND2_X1 _08391_ ( .A1(_01191_ ), .A2(_01202_ ), .ZN(_01203_ ) );
NAND2_X1 _08392_ ( .A1(_01197_ ), .A2(_01198_ ), .ZN(\io_master_araddr [31] ) );
NAND2_X1 _08393_ ( .A1(_01199_ ), .A2(_01200_ ), .ZN(\io_master_araddr [29] ) );
OAI21_X1 _08394_ ( .A(\io_master_araddr [31] ), .B1(\io_master_araddr [30] ), .B2(\io_master_araddr [29] ), .ZN(_01204_ ) );
OAI21_X2 _08395_ ( .A(_01203_ ), .B1(_01196_ ), .B2(_01204_ ), .ZN(_01205_ ) );
NOR3_X1 _08396_ ( .A1(\io_master_araddr [4] ), .A2(\io_master_araddr [5] ), .A3(_01190_ ), .ZN(_01206_ ) );
OR2_X4 _08397_ ( .A1(_01140_ ), .A2(\u_icache.caddr_$_SDFFE_PP0P__Q_29_D_$_MUX__B_A ), .ZN(_01207_ ) );
OAI21_X1 _08398_ ( .A(\u_arbiter.raddr [3] ), .B1(_01138_ ), .B2(\u_arbiter.working ), .ZN(_01208_ ) );
NAND3_X1 _08399_ ( .A1(_01147_ ), .A2(\ca_addr [3] ), .A3(icah_valid ), .ZN(_01209_ ) );
NAND2_X4 _08400_ ( .A1(_01208_ ), .A2(_01209_ ), .ZN(\io_master_araddr [3] ) );
INV_X1 _08401_ ( .A(\u_icache.caddr_$_SDFFE_PP0P__Q_28_D [0] ), .ZN(_01210_ ) );
NAND3_X1 _08402_ ( .A1(_01210_ ), .A2(_00635_ ), .A3(icah_valid ), .ZN(_01211_ ) );
AND3_X2 _08403_ ( .A1(_01207_ ), .A2(\io_master_araddr [3] ), .A3(_01211_ ), .ZN(_01212_ ) );
NOR2_X2 _08404_ ( .A1(_01139_ ), .A2(_01142_ ), .ZN(\io_master_araddr [1] ) );
NOR2_X2 _08405_ ( .A1(\io_master_araddr [1] ), .A2(\io_master_araddr [0] ), .ZN(_01213_ ) );
AND2_X4 _08406_ ( .A1(_01212_ ), .A2(_01213_ ), .ZN(_01214_ ) );
AND3_X2 _08407_ ( .A1(_01206_ ), .A2(_01202_ ), .A3(_01214_ ), .ZN(_01215_ ) );
NAND4_X1 _08408_ ( .A1(_01215_ ), .A2(_01175_ ), .A3(_01160_ ), .A4(_01181_ ), .ZN(_01216_ ) );
NAND4_X1 _08409_ ( .A1(_01146_ ), .A2(_01177_ ), .A3(_01185_ ), .A4(_01150_ ), .ZN(_01217_ ) );
NAND2_X1 _08410_ ( .A1(_01176_ ), .A2(_01180_ ), .ZN(_01218_ ) );
NOR3_X2 _08411_ ( .A1(_01217_ ), .A2(_01159_ ), .A3(_01218_ ), .ZN(_01219_ ) );
OR3_X2 _08412_ ( .A1(\io_master_araddr [4] ), .A2(\io_master_araddr [5] ), .A3(\io_master_araddr [3] ), .ZN(_01220_ ) );
OAI21_X1 _08413_ ( .A(\u_arbiter.raddr [8] ), .B1(_01170_ ), .B2(\u_arbiter.working ), .ZN(_01221_ ) );
NAND3_X1 _08414_ ( .A1(_00635_ ), .A2(\ca_addr [8] ), .A3(icah_valid ), .ZN(_01222_ ) );
NAND4_X1 _08415_ ( .A1(_01220_ ), .A2(\io_master_araddr [6] ), .A3(_01221_ ), .A4(_01222_ ), .ZN(_01223_ ) );
AND3_X2 _08416_ ( .A1(_01219_ ), .A2(_01175_ ), .A3(_01223_ ), .ZN(_01224_ ) );
OAI21_X1 _08417_ ( .A(_01216_ ), .B1(_01224_ ), .B2(_01204_ ), .ZN(_01225_ ) );
INV_X4 _08418_ ( .A(_01225_ ), .ZN(_01226_ ) );
NOR2_X4 _08419_ ( .A1(_01205_ ), .A2(_01226_ ), .ZN(_01227_ ) );
AND2_X4 _08420_ ( .A1(_01227_ ), .A2(\u_lsu.rvalid_clint ), .ZN(_01228_ ) );
INV_X4 _08421_ ( .A(_01228_ ), .ZN(_01229_ ) );
INV_X1 _08422_ ( .A(\u_lsu.u_clint.mtime [47] ), .ZN(_01230_ ) );
INV_X1 _08423_ ( .A(\u_lsu.u_clint.mtime [15] ), .ZN(_01231_ ) );
MUX2_X1 _08424_ ( .A(_01230_ ), .B(_01231_ ), .S(_01214_ ), .Z(_01232_ ) );
OR2_X2 _08425_ ( .A1(_01229_ ), .A2(_01232_ ), .ZN(_01233_ ) );
OAI21_X1 _08426_ ( .A(\io_master_rdata [15] ), .B1(_01205_ ), .B2(_01226_ ), .ZN(_01234_ ) );
AOI21_X1 _08427_ ( .A(_01144_ ), .B1(_01233_ ), .B2(_01234_ ), .ZN(_01235_ ) );
AND2_X2 _08428_ ( .A1(\io_master_araddr [1] ), .A2(\u_arbiter.raddr [0] ), .ZN(_01236_ ) );
INV_X1 _08429_ ( .A(_01236_ ), .ZN(_01237_ ) );
BUF_X8 _08430_ ( .A(_01228_ ), .Z(_01238_ ) );
AND2_X2 _08431_ ( .A1(_01207_ ), .A2(_01211_ ), .ZN(_01239_ ) );
INV_X1 _08432_ ( .A(\u_lsu.u_clint.mtime [31] ), .ZN(_01240_ ) );
NAND4_X1 _08433_ ( .A1(_01239_ ), .A2(_01240_ ), .A3(\io_master_araddr [3] ), .A4(_01213_ ), .ZN(_01241_ ) );
BUF_X4 _08434_ ( .A(_01214_ ), .Z(_01242_ ) );
OAI211_X4 _08435_ ( .A(_01238_ ), .B(_01241_ ), .C1(\u_lsu.u_clint.mtime [63] ), .C2(_01242_ ), .ZN(_01243_ ) );
OAI21_X1 _08436_ ( .A(\io_master_rdata [31] ), .B1(_01205_ ), .B2(_01226_ ), .ZN(_01244_ ) );
AOI21_X2 _08437_ ( .A(_01237_ ), .B1(_01243_ ), .B2(_01244_ ), .ZN(_01245_ ) );
AND2_X1 _08438_ ( .A1(\io_master_araddr [1] ), .A2(_01141_ ), .ZN(_01246_ ) );
INV_X1 _08439_ ( .A(_01246_ ), .ZN(_01247_ ) );
OR2_X1 _08440_ ( .A1(_01242_ ), .A2(\u_lsu.u_clint.mtime [55] ), .ZN(_01248_ ) );
INV_X1 _08441_ ( .A(_01242_ ), .ZN(_01249_ ) );
OAI211_X1 _08442_ ( .A(_01228_ ), .B(_01248_ ), .C1(\u_lsu.u_clint.mtime [23] ), .C2(_01249_ ), .ZN(_01250_ ) );
OAI21_X1 _08443_ ( .A(\io_master_rdata [23] ), .B1(_01205_ ), .B2(_01226_ ), .ZN(_01251_ ) );
AOI21_X1 _08444_ ( .A(_01247_ ), .B1(_01250_ ), .B2(_01251_ ), .ZN(_01252_ ) );
OR3_X4 _08445_ ( .A1(_01235_ ), .A2(_01245_ ), .A3(_01252_ ), .ZN(_01253_ ) );
INV_X2 _08446_ ( .A(_01213_ ), .ZN(_01254_ ) );
OR2_X1 _08447_ ( .A1(_01242_ ), .A2(\u_lsu.u_clint.mtime [39] ), .ZN(_01255_ ) );
OAI211_X1 _08448_ ( .A(_01238_ ), .B(_01255_ ), .C1(\u_lsu.u_clint.mtime [7] ), .C2(_01249_ ), .ZN(_01256_ ) );
OAI21_X1 _08449_ ( .A(\io_master_rdata [7] ), .B1(_01205_ ), .B2(_01226_ ), .ZN(_01257_ ) );
AOI21_X2 _08450_ ( .A(_01254_ ), .B1(_01256_ ), .B2(_01257_ ), .ZN(_01258_ ) );
NOR2_X4 _08451_ ( .A1(_01253_ ), .A2(_01258_ ), .ZN(_01259_ ) );
NOR2_X1 _08452_ ( .A1(_01145_ ), .A2(\u_arbiter.rmask [1] ), .ZN(_01260_ ) );
AND3_X1 _08453_ ( .A1(_01260_ ), .A2(\u_arbiter.rmask [0] ), .A3(\u_arbiter.rsign ), .ZN(_01261_ ) );
INV_X1 _08454_ ( .A(_01261_ ), .ZN(_01262_ ) );
NOR2_X4 _08455_ ( .A1(_01259_ ), .A2(_01262_ ), .ZN(_01263_ ) );
AOI21_X1 _08456_ ( .A(_01144_ ), .B1(_01250_ ), .B2(_01251_ ), .ZN(_01264_ ) );
AOI21_X1 _08457_ ( .A(_01247_ ), .B1(_01243_ ), .B2(_01244_ ), .ZN(_01265_ ) );
CLKBUF_X3 _08458_ ( .A(_01213_ ), .Z(_01266_ ) );
NOR3_X1 _08459_ ( .A1(_01264_ ), .A2(_01265_ ), .A3(_01266_ ), .ZN(_01267_ ) );
AND3_X1 _08460_ ( .A1(_01233_ ), .A2(_01266_ ), .A3(_01234_ ), .ZN(_01268_ ) );
NOR2_X2 _08461_ ( .A1(_01267_ ), .A2(_01268_ ), .ZN(_01269_ ) );
INV_X1 _08462_ ( .A(\u_arbiter.rmask [0] ), .ZN(_01270_ ) );
AND4_X1 _08463_ ( .A1(\u_arbiter.rmask [1] ), .A2(_01149_ ), .A3(_01270_ ), .A4(\u_arbiter.rsign ), .ZN(_01271_ ) );
AND2_X2 _08464_ ( .A1(_01269_ ), .A2(_01271_ ), .ZN(_01272_ ) );
OR2_X4 _08465_ ( .A1(_01263_ ), .A2(_01272_ ), .ZN(_01273_ ) );
BUF_X4 _08466_ ( .A(_01260_ ), .Z(_01274_ ) );
NOR2_X1 _08467_ ( .A1(_01145_ ), .A2(\u_arbiter.rmask [0] ), .ZN(_01275_ ) );
NOR2_X1 _08468_ ( .A1(_01274_ ), .A2(_01275_ ), .ZN(\io_master_arsize [1] ) );
BUF_X4 _08469_ ( .A(_01254_ ), .Z(_01276_ ) );
BUF_X2 _08470_ ( .A(_01276_ ), .Z(_01277_ ) );
AOI21_X1 _08471_ ( .A(_01277_ ), .B1(_01243_ ), .B2(_01244_ ), .ZN(_01278_ ) );
AOI21_X2 _08472_ ( .A(_01273_ ), .B1(\io_master_arsize [1] ), .B2(_01278_ ), .ZN(_01279_ ) );
AOI21_X2 _08473_ ( .A(_01137_ ), .B1(_01279_ ), .B2(fanout_net_9 ), .ZN(\ar_data [31] ) );
MUX2_X1 _08474_ ( .A(io_master_rvalid ), .B(\u_lsu.rvalid_clint ), .S(_01227_ ), .Z(\u_lsu.rvalid ) );
MUX2_X1 _08475_ ( .A(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_A ), .B(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ), .S(_01145_ ), .Z(_01280_ ) );
INV_X1 _08476_ ( .A(fanout_net_9 ), .ZN(_01281_ ) );
NOR2_X1 _08477_ ( .A1(_01280_ ), .A2(_01281_ ), .ZN(_01282_ ) );
NAND3_X2 _08478_ ( .A1(\u_lsu.rvalid ), .A2(\u_lsu.reading ), .A3(_01282_ ), .ZN(_01283_ ) );
NAND4_X1 _08479_ ( .A1(_00760_ ), .A2(_00785_ ), .A3(\u_exu.eopt [0] ), .A4(_00783_ ), .ZN(_01284_ ) );
AND2_X4 _08480_ ( .A1(_01283_ ), .A2(_01284_ ), .ZN(_01285_ ) );
INV_X8 _08481_ ( .A(_01285_ ), .ZN(_01286_ ) );
NAND2_X1 _08482_ ( .A1(_01281_ ), .A2(\ea_ard [2] ), .ZN(_01287_ ) );
NAND2_X1 _08483_ ( .A1(fanout_net_9 ), .A2(\u_arbiter.wbaddr [2] ), .ZN(_01288_ ) );
NAND2_X1 _08484_ ( .A1(_01287_ ), .A2(_01288_ ), .ZN(_01289_ ) );
INV_X1 _08485_ ( .A(_01289_ ), .ZN(_01290_ ) );
XNOR2_X1 _08486_ ( .A(_00948_ ), .B(_01290_ ), .ZN(_01291_ ) );
INV_X2 _08487_ ( .A(_00935_ ), .ZN(_01292_ ) );
NAND2_X1 _08488_ ( .A1(_01281_ ), .A2(\ea_ard [1] ), .ZN(_01293_ ) );
NAND2_X1 _08489_ ( .A1(fanout_net_9 ), .A2(\u_arbiter.wbaddr [1] ), .ZN(_01294_ ) );
NAND2_X1 _08490_ ( .A1(_01293_ ), .A2(_01294_ ), .ZN(_01295_ ) );
INV_X1 _08491_ ( .A(_01295_ ), .ZN(_01296_ ) );
NAND2_X1 _08492_ ( .A1(_01281_ ), .A2(\ea_ard [3] ), .ZN(_01297_ ) );
NAND2_X1 _08493_ ( .A1(\u_arbiter.wbaddr [3] ), .A2(fanout_net_9 ), .ZN(_01298_ ) );
NAND2_X1 _08494_ ( .A1(_01297_ ), .A2(_01298_ ), .ZN(_01299_ ) );
INV_X1 _08495_ ( .A(_01299_ ), .ZN(_01300_ ) );
OAI22_X1 _08496_ ( .A1(_01292_ ), .A2(_01296_ ), .B1(_01043_ ), .B2(_01300_ ), .ZN(_01301_ ) );
NAND2_X1 _08497_ ( .A1(_01281_ ), .A2(\ea_ard [0] ), .ZN(_01302_ ) );
NAND2_X1 _08498_ ( .A1(fanout_net_9 ), .A2(\u_arbiter.wbaddr [0] ), .ZN(_01303_ ) );
NAND2_X1 _08499_ ( .A1(_01302_ ), .A2(_01303_ ), .ZN(_01304_ ) );
INV_X1 _08500_ ( .A(_01304_ ), .ZN(_01305_ ) );
XNOR2_X1 _08501_ ( .A(_00938_ ), .B(_01305_ ), .ZN(_01306_ ) );
BUF_X4 _08502_ ( .A(_00935_ ), .Z(_01307_ ) );
BUF_X2 _08503_ ( .A(_01299_ ), .Z(_01308_ ) );
OAI22_X1 _08504_ ( .A1(_01307_ ), .A2(_01295_ ), .B1(_00944_ ), .B2(_01308_ ), .ZN(_01309_ ) );
NOR4_X1 _08505_ ( .A1(_01291_ ), .A2(_01301_ ), .A3(_01306_ ), .A4(_01309_ ), .ZN(_01310_ ) );
AND2_X4 _08506_ ( .A1(_01286_ ), .A2(_01310_ ), .ZN(_01311_ ) );
INV_X1 _08507_ ( .A(_01311_ ), .ZN(_01312_ ) );
BUF_X4 _08508_ ( .A(_01312_ ), .Z(_01313_ ) );
NOR2_X2 _08509_ ( .A1(\ar_data [31] ), .A2(_01313_ ), .ZN(_01314_ ) );
AND2_X1 _08510_ ( .A1(_00709_ ), .A2(_00737_ ), .ZN(_01315_ ) );
BUF_X4 _08511_ ( .A(_01315_ ), .Z(_01316_ ) );
BUF_X2 _08512_ ( .A(_01316_ ), .Z(_01317_ ) );
BUF_X2 _08513_ ( .A(_01311_ ), .Z(_01318_ ) );
BUF_X4 _08514_ ( .A(_01017_ ), .Z(_01319_ ) );
BUF_X4 _08515_ ( .A(_01319_ ), .Z(_01320_ ) );
BUF_X4 _08516_ ( .A(_00976_ ), .Z(_01321_ ) );
BUF_X4 _08517_ ( .A(_01321_ ), .Z(_01322_ ) );
AOI22_X1 _08518_ ( .A1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01323_ ) );
BUF_X4 _08519_ ( .A(_00948_ ), .Z(_01324_ ) );
BUF_X4 _08520_ ( .A(_01324_ ), .Z(_01325_ ) );
BUF_X4 _08521_ ( .A(_01325_ ), .Z(_01326_ ) );
BUF_X4 _08522_ ( .A(_00965_ ), .Z(_01327_ ) );
BUF_X4 _08523_ ( .A(_01327_ ), .Z(_01328_ ) );
BUF_X4 _08524_ ( .A(_00940_ ), .Z(_01329_ ) );
BUF_X4 _08525_ ( .A(_01329_ ), .Z(_01330_ ) );
BUF_X4 _08526_ ( .A(_01330_ ), .Z(_01331_ ) );
AOI22_X1 _08527_ ( .A1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01332_ ) );
NAND3_X1 _08528_ ( .A1(_01323_ ), .A2(_01326_ ), .A3(_01332_ ), .ZN(_01333_ ) );
BUF_X2 _08529_ ( .A(_00944_ ), .Z(_01334_ ) );
BUF_X4 _08530_ ( .A(_01026_ ), .Z(_01335_ ) );
BUF_X4 _08531_ ( .A(_00938_ ), .Z(_01336_ ) );
BUF_X4 _08532_ ( .A(_01336_ ), .Z(_01337_ ) );
BUF_X4 _08533_ ( .A(_01337_ ), .Z(_01338_ ) );
BUF_X4 _08534_ ( .A(_00933_ ), .Z(_01339_ ) );
BUF_X4 _08535_ ( .A(_00934_ ), .Z(_01340_ ) );
OAI211_X1 _08536_ ( .A(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01338_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_01341_ ) );
BUF_X4 _08537_ ( .A(_00939_ ), .Z(_01342_ ) );
BUF_X4 _08538_ ( .A(_01342_ ), .Z(_01343_ ) );
BUF_X4 _08539_ ( .A(_01307_ ), .Z(_01344_ ) );
BUF_X4 _08540_ ( .A(_01344_ ), .Z(_01345_ ) );
INV_X1 _08541_ ( .A(\u_reg.rf[1][31] ), .ZN(_01346_ ) );
AOI21_X1 _08542_ ( .A(_01343_ ), .B1(_01345_ ), .B2(_01346_ ), .ZN(_01347_ ) );
NOR2_X1 _08543_ ( .A1(_01345_ ), .A2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01348_ ) );
OAI211_X1 _08544_ ( .A(_01335_ ), .B(_01341_ ), .C1(_01347_ ), .C2(_01348_ ), .ZN(_01349_ ) );
NAND3_X1 _08545_ ( .A1(_01333_ ), .A2(_01334_ ), .A3(_01349_ ), .ZN(_01350_ ) );
BUF_X4 _08546_ ( .A(_01319_ ), .Z(_01351_ ) );
BUF_X4 _08547_ ( .A(_01321_ ), .Z(_01352_ ) );
AOI22_X1 _08548_ ( .A1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01353_ ) );
BUF_X4 _08549_ ( .A(_01026_ ), .Z(_01354_ ) );
BUF_X4 _08550_ ( .A(_01330_ ), .Z(_01355_ ) );
AOI22_X1 _08551_ ( .A1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01356_ ) );
NAND3_X1 _08552_ ( .A1(_01353_ ), .A2(_01354_ ), .A3(_01356_ ), .ZN(_01357_ ) );
BUF_X4 _08553_ ( .A(_01319_ ), .Z(_01358_ ) );
BUF_X4 _08554_ ( .A(_01321_ ), .Z(_01359_ ) );
AOI22_X1 _08555_ ( .A1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01360_ ) );
BUF_X4 _08556_ ( .A(_01325_ ), .Z(_01361_ ) );
BUF_X4 _08557_ ( .A(_01327_ ), .Z(_01362_ ) );
BUF_X4 _08558_ ( .A(_01330_ ), .Z(_01363_ ) );
AOI22_X1 _08559_ ( .A1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01364_ ) );
NAND3_X1 _08560_ ( .A1(_01360_ ), .A2(_01361_ ), .A3(_01364_ ), .ZN(_01365_ ) );
BUF_X2 _08561_ ( .A(_01043_ ), .Z(_01366_ ) );
NAND3_X1 _08562_ ( .A1(_01357_ ), .A2(_01365_ ), .A3(_01366_ ), .ZN(_01367_ ) );
AOI21_X1 _08563_ ( .A(_01318_ ), .B1(_01350_ ), .B2(_01367_ ), .ZN(_01368_ ) );
NOR3_X2 _08564_ ( .A1(_01314_ ), .A2(_01317_ ), .A3(_01368_ ), .ZN(_01369_ ) );
BUF_X4 _08565_ ( .A(_00719_ ), .Z(_01370_ ) );
BUF_X2 _08566_ ( .A(_01370_ ), .Z(_01371_ ) );
NAND2_X1 _08567_ ( .A1(_01369_ ), .A2(_01371_ ), .ZN(_01372_ ) );
AND2_X1 _08568_ ( .A1(_00751_ ), .A2(_00757_ ), .ZN(_01373_ ) );
INV_X1 _08569_ ( .A(_01373_ ), .ZN(_01374_ ) );
BUF_X4 _08570_ ( .A(_01374_ ), .Z(_01375_ ) );
AND2_X1 _08571_ ( .A1(_00784_ ), .A2(\u_exu.acsrd [1] ), .ZN(_01376_ ) );
INV_X1 _08572_ ( .A(_01376_ ), .ZN(_01377_ ) );
AND3_X2 _08573_ ( .A1(_00872_ ), .A2(_00639_ ), .A3(_01377_ ), .ZN(_01378_ ) );
INV_X1 _08574_ ( .A(_01378_ ), .ZN(_01379_ ) );
NAND2_X1 _08575_ ( .A1(_01134_ ), .A2(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ), .ZN(_01380_ ) );
AND2_X2 _08576_ ( .A1(_00637_ ), .A2(_01380_ ), .ZN(_01381_ ) );
INV_X1 _08577_ ( .A(_00871_ ), .ZN(_01382_ ) );
OAI21_X1 _08578_ ( .A(_01376_ ), .B1(_01382_ ), .B2(_00978_ ), .ZN(_01383_ ) );
AND2_X1 _08579_ ( .A1(_00784_ ), .A2(\u_exu.acsrd [11] ), .ZN(_01384_ ) );
INV_X1 _08580_ ( .A(_01384_ ), .ZN(_01385_ ) );
NAND3_X1 _08581_ ( .A1(_00639_ ), .A2(\u_idu.imm_auipc_lui [31] ), .A3(_01385_ ), .ZN(_01386_ ) );
AND4_X2 _08582_ ( .A1(_01379_ ), .A2(_01381_ ), .A3(_01383_ ), .A4(_01386_ ), .ZN(_01387_ ) );
NOR2_X1 _08583_ ( .A1(ea_err ), .A2(\u_exu.acsrd [8] ), .ZN(_01388_ ) );
NAND2_X1 _08584_ ( .A1(_01388_ ), .A2(\u_idu.imm_auipc_lui [28] ), .ZN(_01389_ ) );
INV_X1 _08585_ ( .A(\u_exu.acsrd [3] ), .ZN(_01390_ ) );
NOR2_X1 _08586_ ( .A1(_01390_ ), .A2(ea_err ), .ZN(_01391_ ) );
OR3_X1 _08587_ ( .A1(_00638_ ), .A2(_00888_ ), .A3(_01391_ ), .ZN(_01392_ ) );
NAND3_X1 _08588_ ( .A1(_00890_ ), .A2(_00784_ ), .A3(\u_exu.acsrd [2] ), .ZN(_01393_ ) );
NAND2_X1 _08589_ ( .A1(_01392_ ), .A2(_01393_ ), .ZN(_01394_ ) );
NOR3_X1 _08590_ ( .A1(_01390_ ), .A2(\u_idu.imm_auipc_lui [23] ), .A3(ea_err ), .ZN(_01395_ ) );
AND2_X1 _08591_ ( .A1(_00784_ ), .A2(\u_exu.acsrd [2] ), .ZN(_01396_ ) );
AOI21_X1 _08592_ ( .A(_01396_ ), .B1(_00639_ ), .B2(_00890_ ), .ZN(_01397_ ) );
NOR3_X1 _08593_ ( .A1(_01394_ ), .A2(_01395_ ), .A3(_01397_ ), .ZN(_01398_ ) );
AND2_X1 _08594_ ( .A1(_00784_ ), .A2(\u_exu.acsrd [4] ), .ZN(_01399_ ) );
OR3_X1 _08595_ ( .A1(_00638_ ), .A2(_00887_ ), .A3(_01399_ ), .ZN(_01400_ ) );
NAND3_X1 _08596_ ( .A1(_00656_ ), .A2(_00785_ ), .A3(\u_exu.acsrd [5] ), .ZN(_01401_ ) );
NAND3_X1 _08597_ ( .A1(_00887_ ), .A2(_00784_ ), .A3(\u_exu.acsrd [4] ), .ZN(_01402_ ) );
AND3_X1 _08598_ ( .A1(_01400_ ), .A2(_01401_ ), .A3(_01402_ ), .ZN(_01403_ ) );
NAND4_X1 _08599_ ( .A1(_01387_ ), .A2(_01389_ ), .A3(_01398_ ), .A4(_01403_ ), .ZN(_01404_ ) );
NOR2_X1 _08600_ ( .A1(ea_err ), .A2(\u_exu.acsrd [6] ), .ZN(_01405_ ) );
INV_X1 _08601_ ( .A(_01405_ ), .ZN(_01406_ ) );
AOI21_X1 _08602_ ( .A(\u_idu.imm_auipc_lui [26] ), .B1(_00868_ ), .B2(_00757_ ), .ZN(_01407_ ) );
OAI21_X1 _08603_ ( .A(_01406_ ), .B1(_00638_ ), .B2(_01407_ ), .ZN(_01408_ ) );
INV_X1 _08604_ ( .A(\u_exu.acsrd [7] ), .ZN(_01409_ ) );
NOR2_X1 _08605_ ( .A1(_01409_ ), .A2(ea_err ), .ZN(_01410_ ) );
INV_X1 _08606_ ( .A(_01410_ ), .ZN(_01411_ ) );
NAND3_X1 _08607_ ( .A1(_00639_ ), .A2(\u_idu.imm_auipc_lui [27] ), .A3(_01411_ ), .ZN(_01412_ ) );
AND2_X1 _08608_ ( .A1(_00784_ ), .A2(\u_exu.acsrd [5] ), .ZN(_01413_ ) );
INV_X1 _08609_ ( .A(_01413_ ), .ZN(_01414_ ) );
NAND3_X1 _08610_ ( .A1(_00639_ ), .A2(\u_idu.imm_auipc_lui [25] ), .A3(_01414_ ), .ZN(_01415_ ) );
AOI21_X1 _08611_ ( .A(_01406_ ), .B1(_00873_ ), .B2(_00732_ ), .ZN(_01416_ ) );
NOR3_X1 _08612_ ( .A1(_01409_ ), .A2(\u_idu.imm_auipc_lui [27] ), .A3(ea_err ), .ZN(_01417_ ) );
NOR2_X1 _08613_ ( .A1(_01416_ ), .A2(_01417_ ), .ZN(_01418_ ) );
AND4_X1 _08614_ ( .A1(_01408_ ), .A2(_01412_ ), .A3(_01415_ ), .A4(_01418_ ), .ZN(_01419_ ) );
NOR3_X1 _08615_ ( .A1(_00881_ ), .A2(ea_err ), .A3(\u_exu.acsrd [9] ), .ZN(_01420_ ) );
INV_X1 _08616_ ( .A(_01420_ ), .ZN(_01421_ ) );
INV_X1 _08617_ ( .A(_01388_ ), .ZN(_01422_ ) );
NAND3_X1 _08618_ ( .A1(_00640_ ), .A2(_00884_ ), .A3(_01422_ ), .ZN(_01423_ ) );
AND3_X1 _08619_ ( .A1(_01419_ ), .A2(_01421_ ), .A3(_01423_ ), .ZN(_01424_ ) );
AOI22_X1 _08620_ ( .A1(_00637_ ), .A2(ea_err ), .B1(_00868_ ), .B2(_00757_ ), .ZN(_01425_ ) );
AND2_X1 _08621_ ( .A1(_00877_ ), .A2(_01425_ ), .ZN(_01426_ ) );
NOR2_X1 _08622_ ( .A1(ea_err ), .A2(\u_exu.acsrd [0] ), .ZN(_01427_ ) );
XNOR2_X1 _08623_ ( .A(_01426_ ), .B(_01427_ ), .ZN(_01428_ ) );
NAND3_X1 _08624_ ( .A1(_00861_ ), .A2(_00785_ ), .A3(\u_exu.acsrd [10] ), .ZN(_01429_ ) );
NOR2_X1 _08625_ ( .A1(ea_err ), .A2(\u_exu.acsrd [9] ), .ZN(_01430_ ) );
INV_X1 _08626_ ( .A(_01430_ ), .ZN(_01431_ ) );
NAND3_X1 _08627_ ( .A1(_00639_ ), .A2(_00881_ ), .A3(_01431_ ), .ZN(_01432_ ) );
AND2_X1 _08628_ ( .A1(_00784_ ), .A2(\u_exu.acsrd [10] ), .ZN(_01433_ ) );
INV_X1 _08629_ ( .A(_01433_ ), .ZN(_01434_ ) );
NAND3_X1 _08630_ ( .A1(_00639_ ), .A2(\u_idu.imm_auipc_lui [30] ), .A3(_01434_ ), .ZN(_01435_ ) );
NAND3_X1 _08631_ ( .A1(_00662_ ), .A2(_00784_ ), .A3(\u_exu.acsrd [11] ), .ZN(_01436_ ) );
AND4_X1 _08632_ ( .A1(_01429_ ), .A2(_01432_ ), .A3(_01435_ ), .A4(_01436_ ), .ZN(_01437_ ) );
NAND3_X1 _08633_ ( .A1(_01424_ ), .A2(_01428_ ), .A3(_01437_ ), .ZN(_01438_ ) );
OR2_X2 _08634_ ( .A1(_01404_ ), .A2(_01438_ ), .ZN(_01439_ ) );
NOR2_X1 _08635_ ( .A1(_01118_ ), .A2(_01100_ ), .ZN(_01440_ ) );
NOR2_X1 _08636_ ( .A1(_01440_ ), .A2(_00857_ ), .ZN(_01441_ ) );
INV_X1 _08637_ ( .A(_01441_ ), .ZN(_01442_ ) );
BUF_X4 _08638_ ( .A(_01442_ ), .Z(_01443_ ) );
BUF_X4 _08639_ ( .A(_01443_ ), .Z(_01444_ ) );
NOR2_X1 _08640_ ( .A1(_00638_ ), .A2(\u_idu.imm_auipc_lui [22] ), .ZN(_01445_ ) );
INV_X1 _08641_ ( .A(_00869_ ), .ZN(_01446_ ) );
AND4_X1 _08642_ ( .A1(_00732_ ), .A2(_00731_ ), .A3(_00644_ ), .A4(_00752_ ), .ZN(_01447_ ) );
NAND2_X1 _08643_ ( .A1(_01446_ ), .A2(_01447_ ), .ZN(_01448_ ) );
AND2_X1 _08644_ ( .A1(_00640_ ), .A2(_01448_ ), .ZN(_01449_ ) );
AOI211_X1 _08645_ ( .A(_01445_ ), .B(_01449_ ), .C1(\u_idu.imm_auipc_lui [23] ), .C2(_00640_ ), .ZN(_01450_ ) );
BUF_X2 _08646_ ( .A(_01450_ ), .Z(_01451_ ) );
AND2_X1 _08647_ ( .A1(_00872_ ), .A2(_00639_ ), .ZN(_01452_ ) );
NOR2_X1 _08648_ ( .A1(_01452_ ), .A2(_01426_ ), .ZN(_01453_ ) );
BUF_X4 _08649_ ( .A(_01453_ ), .Z(_01454_ ) );
BUF_X2 _08650_ ( .A(_01454_ ), .Z(_01455_ ) );
NAND3_X1 _08651_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][31] ), .A3(_01455_ ), .ZN(_01456_ ) );
NOR4_X1 _08652_ ( .A1(_00872_ ), .A2(\u_idu.imm_auipc_lui [23] ), .A3(\u_idu.imm_auipc_lui [22] ), .A4(_00638_ ), .ZN(_01457_ ) );
CLKBUF_X2 _08653_ ( .A(_01457_ ), .Z(_01458_ ) );
CLKBUF_X2 _08654_ ( .A(_01458_ ), .Z(_01459_ ) );
AND4_X1 _08655_ ( .A1(_00640_ ), .A2(_00877_ ), .A3(_01446_ ), .A4(_01447_ ), .ZN(_01460_ ) );
CLKBUF_X2 _08656_ ( .A(_01460_ ), .Z(_01461_ ) );
CLKBUF_X2 _08657_ ( .A(_01461_ ), .Z(_01462_ ) );
NAND3_X1 _08658_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][31] ), .A3(_01462_ ), .ZN(_01463_ ) );
AND2_X1 _08659_ ( .A1(_01445_ ), .A2(_00888_ ), .ZN(_01464_ ) );
BUF_X4 _08660_ ( .A(_01464_ ), .Z(_01465_ ) );
NOR2_X1 _08661_ ( .A1(_00638_ ), .A2(_01407_ ), .ZN(_01466_ ) );
AND3_X2 _08662_ ( .A1(_01466_ ), .A2(_00731_ ), .A3(_00754_ ), .ZN(_01467_ ) );
NAND4_X1 _08663_ ( .A1(_01454_ ), .A2(\u_csr.csr[2][31] ), .A3(_01465_ ), .A4(_01467_ ), .ZN(_01468_ ) );
NAND3_X1 _08664_ ( .A1(_01456_ ), .A2(_01463_ ), .A3(_01468_ ), .ZN(_01469_ ) );
NAND3_X1 _08665_ ( .A1(_01439_ ), .A2(_01444_ ), .A3(_01469_ ), .ZN(_01470_ ) );
NOR2_X2 _08666_ ( .A1(_01404_ ), .A2(_01438_ ), .ZN(_01471_ ) );
BUF_X4 _08667_ ( .A(_01471_ ), .Z(_01472_ ) );
NAND4_X1 _08668_ ( .A1(_01472_ ), .A2(_00787_ ), .A3(_00786_ ), .A4(_01443_ ), .ZN(_01473_ ) );
AOI21_X1 _08669_ ( .A(_01375_ ), .B1(_01470_ ), .B2(_01473_ ), .ZN(_01474_ ) );
AND2_X1 _08670_ ( .A1(_00742_ ), .A2(_00743_ ), .ZN(_01475_ ) );
NOR2_X1 _08671_ ( .A1(_01475_ ), .A2(_00719_ ), .ZN(_01476_ ) );
AND3_X1 _08672_ ( .A1(_00742_ ), .A2(_00743_ ), .A3(_01374_ ), .ZN(_01477_ ) );
NOR2_X1 _08673_ ( .A1(_01476_ ), .A2(_01477_ ), .ZN(_01478_ ) );
INV_X1 _08674_ ( .A(_01478_ ), .ZN(_01479_ ) );
BUF_X4 _08675_ ( .A(_01479_ ), .Z(_01480_ ) );
AOI221_X4 _08676_ ( .A(_01474_ ), .B1(\de_pc [31] ), .B2(_01480_ ), .C1(_01106_ ), .C2(_01109_ ), .ZN(_01481_ ) );
AND2_X1 _08677_ ( .A1(_00709_ ), .A2(_00898_ ), .ZN(_01482_ ) );
BUF_X4 _08678_ ( .A(_01482_ ), .Z(_01483_ ) );
INV_X2 _08679_ ( .A(_01483_ ), .ZN(_01484_ ) );
BUF_X4 _08680_ ( .A(_01484_ ), .Z(_01485_ ) );
NAND2_X1 _08681_ ( .A1(_01369_ ), .A2(_01485_ ), .ZN(_01486_ ) );
BUF_X4 _08682_ ( .A(_01056_ ), .Z(_01487_ ) );
OR2_X1 _08683_ ( .A1(_00711_ ), .A2(_01075_ ), .ZN(_01488_ ) );
NOR2_X1 _08684_ ( .A1(_01074_ ), .A2(_01488_ ), .ZN(_01489_ ) );
INV_X1 _08685_ ( .A(_01489_ ), .ZN(_01490_ ) );
AND2_X2 _08686_ ( .A1(_01483_ ), .A2(_01490_ ), .ZN(_01491_ ) );
BUF_X4 _08687_ ( .A(_01491_ ), .Z(_01492_ ) );
BUF_X4 _08688_ ( .A(_01489_ ), .Z(_01493_ ) );
AND2_X1 _08689_ ( .A1(_00709_ ), .A2(_01493_ ), .ZN(_01494_ ) );
BUF_X4 _08690_ ( .A(_01494_ ), .Z(_01495_ ) );
NOR2_X1 _08691_ ( .A1(_00692_ ), .A2(_00684_ ), .ZN(_01496_ ) );
AND2_X1 _08692_ ( .A1(_01496_ ), .A2(_00895_ ), .ZN(_01497_ ) );
OR2_X1 _08693_ ( .A1(_01497_ ), .A2(_00860_ ), .ZN(_01498_ ) );
INV_X1 _08694_ ( .A(_01498_ ), .ZN(_01499_ ) );
NAND4_X1 _08695_ ( .A1(_00646_ ), .A2(_00695_ ), .A3(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A4(\u_idu.imm_auipc_lui [31] ), .ZN(_01500_ ) );
NOR2_X1 _08696_ ( .A1(_00899_ ), .A2(_01500_ ), .ZN(_01501_ ) );
INV_X1 _08697_ ( .A(_01501_ ), .ZN(_01502_ ) );
OR3_X1 _08698_ ( .A1(_00693_ ), .A2(_00860_ ), .A3(_01084_ ), .ZN(_01503_ ) );
OAI221_X1 _08699_ ( .A(_01502_ ), .B1(_00860_ ), .B2(_00900_ ), .C1(_00898_ ), .C2(_01503_ ), .ZN(_01504_ ) );
OR2_X1 _08700_ ( .A1(_01499_ ), .A2(_01504_ ), .ZN(_01505_ ) );
AOI221_X1 _08701_ ( .A(_01487_ ), .B1(\de_pc [31] ), .B2(_01492_ ), .C1(_01495_ ), .C2(_01505_ ), .ZN(_01506_ ) );
AOI221_X1 _08702_ ( .A(_00893_ ), .B1(_01372_ ), .B2(_01481_ ), .C1(_01486_ ), .C2(_01506_ ), .ZN(_00129_ ) );
INV_X1 _08703_ ( .A(_01492_ ), .ZN(_01507_ ) );
INV_X1 _08704_ ( .A(\de_pc [30] ), .ZN(_01508_ ) );
INV_X1 _08705_ ( .A(_01494_ ), .ZN(_01509_ ) );
CLKBUF_X2 _08706_ ( .A(_01498_ ), .Z(_01510_ ) );
BUF_X4 _08707_ ( .A(_00713_ ), .Z(_01511_ ) );
BUF_X4 _08708_ ( .A(_00714_ ), .Z(_01512_ ) );
NAND3_X1 _08709_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [30] ), .A3(_01512_ ), .ZN(_01513_ ) );
AOI21_X1 _08710_ ( .A(_00719_ ), .B1(_00711_ ), .B2(_01094_ ), .ZN(_01514_ ) );
NOR2_X1 _08711_ ( .A1(_01514_ ), .A2(_00860_ ), .ZN(_01515_ ) );
INV_X1 _08712_ ( .A(_01515_ ), .ZN(_01516_ ) );
CLKBUF_X2 _08713_ ( .A(_01516_ ), .Z(_01517_ ) );
AND3_X1 _08714_ ( .A1(_01510_ ), .A2(_01513_ ), .A3(_01517_ ), .ZN(_01518_ ) );
OAI22_X1 _08715_ ( .A1(_01507_ ), .A2(_01508_ ), .B1(_01509_ ), .B2(_01518_ ), .ZN(_01519_ ) );
AND3_X1 _08716_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [30] ), .ZN(_01520_ ) );
BUF_X4 _08717_ ( .A(_01135_ ), .Z(_01521_ ) );
AOI211_X1 _08718_ ( .A(fanout_net_9 ), .B(_01520_ ), .C1(\ea_addr [30] ), .C2(_01521_ ), .ZN(_01522_ ) );
BUF_X16 _08719_ ( .A(_01273_ ), .Z(_01523_ ) );
BUF_X2 _08720_ ( .A(_01266_ ), .Z(_01524_ ) );
AND2_X2 _08721_ ( .A1(_01524_ ), .A2(\io_master_arsize [1] ), .ZN(_01525_ ) );
BUF_X4 _08722_ ( .A(_01227_ ), .Z(_01526_ ) );
BUF_X8 _08723_ ( .A(_01526_ ), .Z(_01527_ ) );
OR2_X1 _08724_ ( .A1(_01527_ ), .A2(\io_master_rdata [30] ), .ZN(_01528_ ) );
BUF_X2 _08725_ ( .A(_01242_ ), .Z(_01529_ ) );
MUX2_X1 _08726_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ), .B(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_31_A_$_ANDNOT__Y_B ), .S(_01529_ ), .Z(_01530_ ) );
OAI21_X1 _08727_ ( .A(_01527_ ), .B1(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .B2(_01530_ ), .ZN(_01531_ ) );
AND2_X4 _08728_ ( .A1(_01528_ ), .A2(_01531_ ), .ZN(_01532_ ) );
AOI21_X4 _08729_ ( .A(_01523_ ), .B1(_01525_ ), .B2(_01532_ ), .ZN(_01533_ ) );
AOI21_X4 _08730_ ( .A(_01522_ ), .B1(_01533_ ), .B2(fanout_net_9 ), .ZN(\ar_data [30] ) );
OR2_X2 _08731_ ( .A1(\ar_data [30] ), .A2(_01313_ ), .ZN(_01534_ ) );
INV_X1 _08732_ ( .A(_01316_ ), .ZN(_01535_ ) );
BUF_X2 _08733_ ( .A(_01312_ ), .Z(_01536_ ) );
BUF_X4 _08734_ ( .A(_01319_ ), .Z(_01537_ ) );
BUF_X4 _08735_ ( .A(_01321_ ), .Z(_01538_ ) );
AOI22_X1 _08736_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01539_ ) );
BUF_X4 _08737_ ( .A(_00965_ ), .Z(_01540_ ) );
BUF_X4 _08738_ ( .A(_01540_ ), .Z(_01541_ ) );
BUF_X4 _08739_ ( .A(_01330_ ), .Z(_01542_ ) );
AOI22_X1 _08740_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01543_ ) );
NAND3_X1 _08741_ ( .A1(_01539_ ), .A2(_01326_ ), .A3(_01543_ ), .ZN(_01544_ ) );
BUF_X4 _08742_ ( .A(_01292_ ), .Z(_01545_ ) );
BUF_X4 _08743_ ( .A(_01545_ ), .Z(_01546_ ) );
BUF_X4 _08744_ ( .A(_01337_ ), .Z(_01547_ ) );
NAND3_X1 _08745_ ( .A1(_01546_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01547_ ), .ZN(_01548_ ) );
BUF_X4 _08746_ ( .A(_01344_ ), .Z(_01549_ ) );
NOR2_X1 _08747_ ( .A1(_01549_ ), .A2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01550_ ) );
BUF_X4 _08748_ ( .A(_01344_ ), .Z(_01551_ ) );
INV_X1 _08749_ ( .A(\u_reg.rf[1][30] ), .ZN(_01552_ ) );
AOI21_X1 _08750_ ( .A(_01343_ ), .B1(_01551_ ), .B2(_01552_ ), .ZN(_01553_ ) );
OAI211_X1 _08751_ ( .A(_01548_ ), .B(_01354_ ), .C1(_01550_ ), .C2(_01553_ ), .ZN(_01554_ ) );
AND3_X1 _08752_ ( .A1(_01544_ ), .A2(_01334_ ), .A3(_01554_ ), .ZN(_01555_ ) );
AOI22_X1 _08753_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01556_ ) );
BUF_X4 _08754_ ( .A(_01026_ ), .Z(_01557_ ) );
BUF_X4 _08755_ ( .A(_01557_ ), .Z(_01558_ ) );
BUF_X4 _08756_ ( .A(_01327_ ), .Z(_01559_ ) );
AOI22_X1 _08757_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01560_ ) );
NAND3_X1 _08758_ ( .A1(_01556_ ), .A2(_01558_ ), .A3(_01560_ ), .ZN(_01561_ ) );
AOI22_X1 _08759_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01562_ ) );
AOI22_X1 _08760_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01563_ ) );
NAND3_X1 _08761_ ( .A1(_01562_ ), .A2(_01326_ ), .A3(_01563_ ), .ZN(_01564_ ) );
AND3_X1 _08762_ ( .A1(_01561_ ), .A2(_01564_ ), .A3(_01366_ ), .ZN(_01565_ ) );
OAI21_X1 _08763_ ( .A(_01536_ ), .B1(_01555_ ), .B2(_01565_ ), .ZN(_01566_ ) );
AND3_X2 _08764_ ( .A1(_01534_ ), .A2(_01535_ ), .A3(_01566_ ), .ZN(_01567_ ) );
AOI21_X1 _08765_ ( .A(_01519_ ), .B1(_01567_ ), .B2(_01485_ ), .ZN(_01568_ ) );
AND2_X2 _08766_ ( .A1(_01055_ ), .A2(_00891_ ), .ZN(_01569_ ) );
INV_X1 _08767_ ( .A(_01569_ ), .ZN(_01570_ ) );
NOR2_X1 _08768_ ( .A1(_01568_ ), .A2(_01570_ ), .ZN(_01571_ ) );
INV_X1 _08769_ ( .A(_01069_ ), .ZN(_01572_ ) );
NAND2_X1 _08770_ ( .A1(_01567_ ), .A2(_01371_ ), .ZN(_01573_ ) );
NOR2_X1 _08771_ ( .A1(_01471_ ), .A2(_01441_ ), .ZN(_01574_ ) );
BUF_X4 _08772_ ( .A(_01574_ ), .Z(_01575_ ) );
BUF_X4 _08773_ ( .A(_01575_ ), .Z(_01576_ ) );
BUF_X4 _08774_ ( .A(_01450_ ), .Z(_01577_ ) );
BUF_X2 _08775_ ( .A(_01577_ ), .Z(_01578_ ) );
BUF_X2 _08776_ ( .A(_01455_ ), .Z(_01579_ ) );
AND3_X1 _08777_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][30] ), .A3(_01579_ ), .ZN(_01580_ ) );
AND3_X1 _08778_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][30] ), .A3(_01462_ ), .ZN(_01581_ ) );
AND2_X2 _08779_ ( .A1(_01453_ ), .A2(_01464_ ), .ZN(_01582_ ) );
BUF_X4 _08780_ ( .A(_01582_ ), .Z(_01583_ ) );
BUF_X4 _08781_ ( .A(_01583_ ), .Z(_01584_ ) );
NAND4_X1 _08782_ ( .A1(_00656_ ), .A2(_00886_ ), .A3(\u_idu.imm_auipc_lui [28] ), .A4(\u_idu.imm_auipc_lui [29] ), .ZN(_01585_ ) );
NOR4_X1 _08783_ ( .A1(_01585_ ), .A2(_00662_ ), .A3(_00887_ ), .A4(_00861_ ), .ZN(_01586_ ) );
AND3_X2 _08784_ ( .A1(_00640_ ), .A2(_01407_ ), .A3(_01586_ ), .ZN(_01587_ ) );
BUF_X4 _08785_ ( .A(_01587_ ), .Z(_01588_ ) );
AOI21_X1 _08786_ ( .A(_01581_ ), .B1(_01584_ ), .B2(_01588_ ), .ZN(_01589_ ) );
BUF_X4 _08787_ ( .A(_00754_ ), .Z(_01590_ ) );
AND2_X2 _08788_ ( .A1(_01466_ ), .A2(_00731_ ), .ZN(_01591_ ) );
BUF_X2 _08789_ ( .A(_01591_ ), .Z(_01592_ ) );
NAND4_X1 _08790_ ( .A1(_01584_ ), .A2(\u_csr.csr[2][30] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_01593_ ) );
NAND2_X1 _08791_ ( .A1(_01589_ ), .A2(_01593_ ), .ZN(_01594_ ) );
OAI21_X1 _08792_ ( .A(_01576_ ), .B1(_01580_ ), .B2(_01594_ ), .ZN(_01595_ ) );
BUF_X2 _08793_ ( .A(_01472_ ), .Z(_01596_ ) );
BUF_X2 _08794_ ( .A(_01444_ ), .Z(_01597_ ) );
NAND4_X1 _08795_ ( .A1(_01596_ ), .A2(_00791_ ), .A3(_00790_ ), .A4(_01597_ ), .ZN(_01598_ ) );
AOI21_X1 _08796_ ( .A(_01375_ ), .B1(_01595_ ), .B2(_01598_ ), .ZN(_01599_ ) );
AOI21_X1 _08797_ ( .A(_01599_ ), .B1(\de_pc [30] ), .B2(_01480_ ), .ZN(_01600_ ) );
AOI21_X1 _08798_ ( .A(_01572_ ), .B1(_01573_ ), .B2(_01600_ ), .ZN(_01601_ ) );
OR2_X1 _08799_ ( .A1(_01571_ ), .A2(_01601_ ), .ZN(_00130_ ) );
AND3_X1 _08800_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [21] ), .ZN(_01602_ ) );
AOI211_X1 _08801_ ( .A(fanout_net_9 ), .B(_01602_ ), .C1(\ea_addr [21] ), .C2(_01136_ ), .ZN(_01603_ ) );
BUF_X8 _08802_ ( .A(_01263_ ), .Z(_01604_ ) );
OR2_X1 _08803_ ( .A1(_01529_ ), .A2(\u_lsu.u_clint.mtime [53] ), .ZN(_01605_ ) );
OAI211_X1 _08804_ ( .A(_01238_ ), .B(_01605_ ), .C1(\u_lsu.u_clint.mtime [21] ), .C2(_01249_ ), .ZN(_01606_ ) );
BUF_X2 _08805_ ( .A(_01205_ ), .Z(_01607_ ) );
BUF_X2 _08806_ ( .A(_01226_ ), .Z(_01608_ ) );
OAI21_X1 _08807_ ( .A(\io_master_rdata [21] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_01609_ ) );
AND2_X1 _08808_ ( .A1(_01606_ ), .A2(_01609_ ), .ZN(_01610_ ) );
OR2_X1 _08809_ ( .A1(_01529_ ), .A2(\u_lsu.u_clint.mtime [61] ), .ZN(_01611_ ) );
OAI211_X1 _08810_ ( .A(_01238_ ), .B(_01611_ ), .C1(\u_lsu.u_clint.mtime [29] ), .C2(_01249_ ), .ZN(_01612_ ) );
OAI21_X1 _08811_ ( .A(\io_master_rdata [29] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_01613_ ) );
NAND2_X2 _08812_ ( .A1(_01612_ ), .A2(_01613_ ), .ZN(_01614_ ) );
NAND2_X1 _08813_ ( .A1(_01614_ ), .A2(_01143_ ), .ZN(_01615_ ) );
MUX2_X2 _08814_ ( .A(_01610_ ), .B(_01615_ ), .S(_01254_ ), .Z(_01616_ ) );
NOR3_X1 _08815_ ( .A1(_01616_ ), .A2(_01274_ ), .A3(_01275_ ), .ZN(_01617_ ) );
NOR3_X1 _08816_ ( .A1(_01604_ ), .A2(_01272_ ), .A3(_01617_ ), .ZN(_01618_ ) );
AOI21_X2 _08817_ ( .A(_01603_ ), .B1(_01618_ ), .B2(fanout_net_9 ), .ZN(\ar_data [21] ) );
NOR2_X1 _08818_ ( .A1(\ar_data [21] ), .A2(_01313_ ), .ZN(_01619_ ) );
AOI22_X1 _08819_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01620_ ) );
AOI22_X1 _08820_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01621_ ) );
NAND3_X1 _08821_ ( .A1(_01620_ ), .A2(_01326_ ), .A3(_01621_ ), .ZN(_01622_ ) );
OAI211_X1 _08822_ ( .A(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01338_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_01623_ ) );
INV_X1 _08823_ ( .A(\u_reg.rf[1][21] ), .ZN(_01624_ ) );
AOI21_X1 _08824_ ( .A(_01343_ ), .B1(_01345_ ), .B2(_01624_ ), .ZN(_01625_ ) );
NOR2_X1 _08825_ ( .A1(_01345_ ), .A2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01626_ ) );
OAI211_X1 _08826_ ( .A(_01335_ ), .B(_01623_ ), .C1(_01625_ ), .C2(_01626_ ), .ZN(_01627_ ) );
NAND3_X1 _08827_ ( .A1(_01622_ ), .A2(_01334_ ), .A3(_01627_ ), .ZN(_01628_ ) );
AOI22_X1 _08828_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01629_ ) );
AOI22_X1 _08829_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01630_ ) );
NAND3_X1 _08830_ ( .A1(_01629_ ), .A2(_01354_ ), .A3(_01630_ ), .ZN(_01631_ ) );
AOI22_X1 _08831_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01632_ ) );
BUF_X4 _08832_ ( .A(_01324_ ), .Z(_01633_ ) );
BUF_X4 _08833_ ( .A(_01327_ ), .Z(_01634_ ) );
AOI22_X1 _08834_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01635_ ) );
NAND3_X1 _08835_ ( .A1(_01632_ ), .A2(_01633_ ), .A3(_01635_ ), .ZN(_01636_ ) );
NAND3_X1 _08836_ ( .A1(_01631_ ), .A2(_01636_ ), .A3(_01366_ ), .ZN(_01637_ ) );
AOI21_X1 _08837_ ( .A(_01318_ ), .B1(_01628_ ), .B2(_01637_ ), .ZN(_01638_ ) );
NOR3_X2 _08838_ ( .A1(_01619_ ), .A2(_01317_ ), .A3(_01638_ ), .ZN(_01639_ ) );
NAND2_X1 _08839_ ( .A1(_01639_ ), .A2(_01371_ ), .ZN(_01640_ ) );
AND2_X1 _08840_ ( .A1(_01582_ ), .A2(_01587_ ), .ZN(_01641_ ) );
INV_X1 _08841_ ( .A(_01464_ ), .ZN(_01642_ ) );
NAND4_X1 _08842_ ( .A1(_00872_ ), .A2(_00639_ ), .A3(_00873_ ), .A4(_00877_ ), .ZN(_01643_ ) );
NOR2_X1 _08843_ ( .A1(_01642_ ), .A2(_01643_ ), .ZN(_01644_ ) );
AND2_X1 _08844_ ( .A1(_01644_ ), .A2(_01587_ ), .ZN(_01645_ ) );
NOR2_X1 _08845_ ( .A1(_01641_ ), .A2(_01645_ ), .ZN(_01646_ ) );
BUF_X2 _08846_ ( .A(_01454_ ), .Z(_01647_ ) );
BUF_X4 _08847_ ( .A(_01465_ ), .Z(_01648_ ) );
BUF_X4 _08848_ ( .A(_01467_ ), .Z(_01649_ ) );
NAND4_X1 _08849_ ( .A1(_01647_ ), .A2(\u_csr.csr[2][21] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_01650_ ) );
BUF_X4 _08850_ ( .A(_01454_ ), .Z(_01651_ ) );
NAND3_X1 _08851_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][21] ), .A3(_01651_ ), .ZN(_01652_ ) );
BUF_X2 _08852_ ( .A(_01465_ ), .Z(_01653_ ) );
BUF_X2 _08853_ ( .A(_01426_ ), .Z(_01654_ ) );
AOI22_X2 _08854_ ( .A1(_00640_ ), .A2(_01448_ ), .B1(fanout_net_20 ), .B2(_00871_ ), .ZN(_01655_ ) );
NAND4_X1 _08855_ ( .A1(_01653_ ), .A2(\u_csr.csr[0][21] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_01656_ ) );
NAND4_X1 _08856_ ( .A1(_01646_ ), .A2(_01650_ ), .A3(_01652_ ), .A4(_01656_ ), .ZN(_01657_ ) );
NAND2_X1 _08857_ ( .A1(_01575_ ), .A2(_01657_ ), .ZN(_01658_ ) );
NAND4_X1 _08858_ ( .A1(_01472_ ), .A2(_00793_ ), .A3(_00792_ ), .A4(_01443_ ), .ZN(_01659_ ) );
AOI21_X1 _08859_ ( .A(_01375_ ), .B1(_01658_ ), .B2(_01659_ ), .ZN(_01660_ ) );
AOI221_X4 _08860_ ( .A(_01660_ ), .B1(\de_pc [21] ), .B2(_01480_ ), .C1(_01106_ ), .C2(_01109_ ), .ZN(_01661_ ) );
NAND2_X1 _08861_ ( .A1(_01639_ ), .A2(_01485_ ), .ZN(_01662_ ) );
NAND3_X1 _08862_ ( .A1(_01511_ ), .A2(fanout_net_20 ), .A3(_01512_ ), .ZN(_01663_ ) );
NAND3_X1 _08863_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_01663_ ), .ZN(_01664_ ) );
AOI221_X1 _08864_ ( .A(_01487_ ), .B1(\de_pc [21] ), .B2(_01492_ ), .C1(_01495_ ), .C2(_01664_ ), .ZN(_01665_ ) );
AOI221_X1 _08865_ ( .A(_00893_ ), .B1(_01640_ ), .B2(_01661_ ), .C1(_01662_ ), .C2(_01665_ ), .ZN(_00131_ ) );
AND3_X1 _08866_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [20] ), .ZN(_01666_ ) );
AOI211_X1 _08867_ ( .A(fanout_net_9 ), .B(_01666_ ), .C1(\ea_addr [20] ), .C2(_01521_ ), .ZN(_01667_ ) );
OR2_X1 _08868_ ( .A1(_01526_ ), .A2(\io_master_rdata [28] ), .ZN(_01668_ ) );
CLKBUF_X2 _08869_ ( .A(_01212_ ), .Z(_01669_ ) );
AND3_X1 _08870_ ( .A1(_01669_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ), .A3(_01266_ ), .ZN(_01670_ ) );
INV_X1 _08871_ ( .A(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .ZN(_01671_ ) );
INV_X1 _08872_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ), .ZN(_01672_ ) );
OAI21_X1 _08873_ ( .A(_01671_ ), .B1(_01529_ ), .B2(_01672_ ), .ZN(_01673_ ) );
OAI21_X1 _08874_ ( .A(_01527_ ), .B1(_01670_ ), .B2(_01673_ ), .ZN(_01674_ ) );
AND2_X1 _08875_ ( .A1(_01668_ ), .A2(_01674_ ), .ZN(_01675_ ) );
INV_X1 _08876_ ( .A(\io_master_araddr [0] ), .ZN(_01676_ ) );
OR2_X1 _08877_ ( .A1(_01675_ ), .A2(_01676_ ), .ZN(_01677_ ) );
OR2_X1 _08878_ ( .A1(_01526_ ), .A2(\io_master_rdata [20] ), .ZN(_01678_ ) );
AND3_X1 _08879_ ( .A1(_01669_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ), .A3(_01266_ ), .ZN(_01679_ ) );
INV_X1 _08880_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_10_A_$_ANDNOT__Y_B ), .ZN(_01680_ ) );
OAI21_X1 _08881_ ( .A(_01671_ ), .B1(_01529_ ), .B2(_01680_ ), .ZN(_01681_ ) );
OAI21_X1 _08882_ ( .A(_01526_ ), .B1(_01679_ ), .B2(_01681_ ), .ZN(_01682_ ) );
AOI21_X1 _08883_ ( .A(_01276_ ), .B1(_01678_ ), .B2(_01682_ ), .ZN(_01683_ ) );
NOR4_X1 _08884_ ( .A1(_01683_ ), .A2(\io_master_araddr [1] ), .A3(_01274_ ), .A4(_01275_ ), .ZN(_01684_ ) );
AOI21_X4 _08885_ ( .A(_01523_ ), .B1(_01677_ ), .B2(_01684_ ), .ZN(_01685_ ) );
AOI21_X4 _08886_ ( .A(_01667_ ), .B1(_01685_ ), .B2(fanout_net_9 ), .ZN(\ar_data [20] ) );
BUF_X4 _08887_ ( .A(_01312_ ), .Z(_01686_ ) );
NOR2_X2 _08888_ ( .A1(\ar_data [20] ), .A2(_01686_ ), .ZN(_01687_ ) );
BUF_X4 _08889_ ( .A(_01311_ ), .Z(_01688_ ) );
AOI22_X1 _08890_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01689_ ) );
AOI22_X1 _08891_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01690_ ) );
NAND3_X1 _08892_ ( .A1(_01689_ ), .A2(_01326_ ), .A3(_01690_ ), .ZN(_01691_ ) );
NAND3_X1 _08893_ ( .A1(_01546_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01338_ ), .ZN(_01692_ ) );
NOR2_X1 _08894_ ( .A1(_01551_ ), .A2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01693_ ) );
BUF_X4 _08895_ ( .A(_01342_ ), .Z(_01694_ ) );
INV_X1 _08896_ ( .A(\u_reg.rf[1][20] ), .ZN(_01695_ ) );
AOI21_X1 _08897_ ( .A(_01694_ ), .B1(_01345_ ), .B2(_01695_ ), .ZN(_01696_ ) );
OAI211_X1 _08898_ ( .A(_01692_ ), .B(_01335_ ), .C1(_01693_ ), .C2(_01696_ ), .ZN(_01697_ ) );
NAND3_X1 _08899_ ( .A1(_01691_ ), .A2(_01334_ ), .A3(_01697_ ), .ZN(_01698_ ) );
AOI22_X1 _08900_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01699_ ) );
AOI22_X1 _08901_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01700_ ) );
NAND3_X1 _08902_ ( .A1(_01699_ ), .A2(_01354_ ), .A3(_01700_ ), .ZN(_01701_ ) );
AOI22_X1 _08903_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01702_ ) );
AOI22_X1 _08904_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01703_ ) );
NAND3_X1 _08905_ ( .A1(_01702_ ), .A2(_01633_ ), .A3(_01703_ ), .ZN(_01704_ ) );
BUF_X2 _08906_ ( .A(_01043_ ), .Z(_01705_ ) );
NAND3_X1 _08907_ ( .A1(_01701_ ), .A2(_01704_ ), .A3(_01705_ ), .ZN(_01706_ ) );
AOI21_X1 _08908_ ( .A(_01688_ ), .B1(_01698_ ), .B2(_01706_ ), .ZN(_01707_ ) );
NOR3_X2 _08909_ ( .A1(_01687_ ), .A2(_01317_ ), .A3(_01707_ ), .ZN(_01708_ ) );
NAND2_X1 _08910_ ( .A1(_01708_ ), .A2(_01371_ ), .ZN(_01709_ ) );
NAND4_X1 _08911_ ( .A1(_01455_ ), .A2(\u_csr.csr[2][20] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_01710_ ) );
NAND3_X1 _08912_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][20] ), .A3(_01647_ ), .ZN(_01711_ ) );
NAND4_X1 _08913_ ( .A1(_01653_ ), .A2(\u_csr.csr[0][20] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_01712_ ) );
NAND4_X1 _08914_ ( .A1(_01646_ ), .A2(_01710_ ), .A3(_01711_ ), .A4(_01712_ ), .ZN(_01713_ ) );
NAND2_X1 _08915_ ( .A1(_01576_ ), .A2(_01713_ ), .ZN(_01714_ ) );
BUF_X4 _08916_ ( .A(_01442_ ), .Z(_01715_ ) );
NAND4_X1 _08917_ ( .A1(_01596_ ), .A2(_00795_ ), .A3(_00794_ ), .A4(_01715_ ), .ZN(_01716_ ) );
AOI21_X1 _08918_ ( .A(_01375_ ), .B1(_01714_ ), .B2(_01716_ ), .ZN(_01717_ ) );
AOI221_X4 _08919_ ( .A(_01717_ ), .B1(\de_pc [20] ), .B2(_01480_ ), .C1(_01106_ ), .C2(_01109_ ), .ZN(_01718_ ) );
NAND2_X1 _08920_ ( .A1(_01708_ ), .A2(_01485_ ), .ZN(_01719_ ) );
BUF_X2 _08921_ ( .A(_01494_ ), .Z(_01720_ ) );
NAND3_X1 _08922_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(_01512_ ), .ZN(_01721_ ) );
NAND3_X1 _08923_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_01721_ ), .ZN(_01722_ ) );
AOI221_X1 _08924_ ( .A(_01487_ ), .B1(\de_pc [20] ), .B2(_01492_ ), .C1(_01720_ ), .C2(_01722_ ), .ZN(_01723_ ) );
AOI221_X1 _08925_ ( .A(_00893_ ), .B1(_01709_ ), .B2(_01718_ ), .C1(_01719_ ), .C2(_01723_ ), .ZN(_00132_ ) );
AND3_X1 _08926_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [19] ), .ZN(_01724_ ) );
AOI211_X1 _08927_ ( .A(fanout_net_9 ), .B(_01724_ ), .C1(\ea_addr [19] ), .C2(_01136_ ), .ZN(_01725_ ) );
INV_X1 _08928_ ( .A(\u_lsu.u_clint.mtime [19] ), .ZN(_01726_ ) );
NAND4_X1 _08929_ ( .A1(_01239_ ), .A2(_01726_ ), .A3(\io_master_araddr [3] ), .A4(_01213_ ), .ZN(_01727_ ) );
OAI211_X1 _08930_ ( .A(_01238_ ), .B(_01727_ ), .C1(\u_lsu.u_clint.mtime [51] ), .C2(_01529_ ), .ZN(_01728_ ) );
OAI21_X1 _08931_ ( .A(\io_master_rdata [19] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_01729_ ) );
AND2_X1 _08932_ ( .A1(_01728_ ), .A2(_01729_ ), .ZN(_01730_ ) );
INV_X1 _08933_ ( .A(\u_lsu.u_clint.mtime [27] ), .ZN(_01731_ ) );
NAND4_X1 _08934_ ( .A1(_01239_ ), .A2(_01731_ ), .A3(\io_master_araddr [3] ), .A4(_01266_ ), .ZN(_01732_ ) );
BUF_X4 _08935_ ( .A(_01242_ ), .Z(_01733_ ) );
OAI211_X2 _08936_ ( .A(_01238_ ), .B(_01732_ ), .C1(\u_lsu.u_clint.mtime [59] ), .C2(_01733_ ), .ZN(_01734_ ) );
OAI21_X1 _08937_ ( .A(\io_master_rdata [27] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_01735_ ) );
NAND2_X2 _08938_ ( .A1(_01734_ ), .A2(_01735_ ), .ZN(_01736_ ) );
NAND2_X1 _08939_ ( .A1(_01736_ ), .A2(_01143_ ), .ZN(_01737_ ) );
MUX2_X1 _08940_ ( .A(_01730_ ), .B(_01737_ ), .S(_01254_ ), .Z(_01738_ ) );
NOR3_X1 _08941_ ( .A1(_01738_ ), .A2(_01274_ ), .A3(_01275_ ), .ZN(_01739_ ) );
NOR3_X1 _08942_ ( .A1(_01604_ ), .A2(_01272_ ), .A3(_01739_ ), .ZN(_01740_ ) );
AOI21_X2 _08943_ ( .A(_01725_ ), .B1(_01740_ ), .B2(fanout_net_9 ), .ZN(\ar_data [19] ) );
NOR2_X1 _08944_ ( .A1(\ar_data [19] ), .A2(_01686_ ), .ZN(_01741_ ) );
AOI22_X1 _08945_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01017_ ), .B1(_01321_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01742_ ) );
AOI22_X1 _08946_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01327_ ), .B1(_01329_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01743_ ) );
AND3_X1 _08947_ ( .A1(_01742_ ), .A2(_01324_ ), .A3(_01743_ ), .ZN(_01744_ ) );
OAI21_X1 _08948_ ( .A(_01336_ ), .B1(_01292_ ), .B2(\u_reg.rf[1][19] ), .ZN(_01745_ ) );
OR2_X1 _08949_ ( .A1(_01307_ ), .A2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01746_ ) );
AOI221_X4 _08950_ ( .A(_01324_ ), .B1(_01329_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(_01745_ ), .C2(_01746_ ), .ZN(_01747_ ) );
OR3_X1 _08951_ ( .A1(_01744_ ), .A2(_01043_ ), .A3(_01747_ ), .ZN(_01748_ ) );
BUF_X4 _08952_ ( .A(_01017_ ), .Z(_01749_ ) );
BUF_X4 _08953_ ( .A(_00976_ ), .Z(_01750_ ) );
AOI22_X1 _08954_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01751_ ) );
BUF_X4 _08955_ ( .A(_00965_ ), .Z(_01752_ ) );
BUF_X4 _08956_ ( .A(_01329_ ), .Z(_01753_ ) );
AOI22_X1 _08957_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01752_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01754_ ) );
AOI21_X1 _08958_ ( .A(_01557_ ), .B1(_01751_ ), .B2(_01754_ ), .ZN(_01755_ ) );
BUF_X2 _08959_ ( .A(_01324_ ), .Z(_01756_ ) );
BUF_X4 _08960_ ( .A(_01017_ ), .Z(_01757_ ) );
BUF_X4 _08961_ ( .A(_00976_ ), .Z(_01758_ ) );
AOI22_X1 _08962_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01759_ ) );
BUF_X4 _08963_ ( .A(_01329_ ), .Z(_01760_ ) );
AOI22_X1 _08964_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01752_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01761_ ) );
AOI21_X1 _08965_ ( .A(_01756_ ), .B1(_01759_ ), .B2(_01761_ ), .ZN(_01762_ ) );
OAI21_X1 _08966_ ( .A(_01366_ ), .B1(_01755_ ), .B2(_01762_ ), .ZN(_01763_ ) );
AOI21_X1 _08967_ ( .A(_01688_ ), .B1(_01748_ ), .B2(_01763_ ), .ZN(_01764_ ) );
NOR3_X2 _08968_ ( .A1(_01741_ ), .A2(_01317_ ), .A3(_01764_ ), .ZN(_01765_ ) );
NAND2_X1 _08969_ ( .A1(_01765_ ), .A2(_01371_ ), .ZN(_01766_ ) );
BUF_X4 _08970_ ( .A(_01374_ ), .Z(_01767_ ) );
AND3_X1 _08971_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][19] ), .A3(_01461_ ), .ZN(_01768_ ) );
AOI21_X1 _08972_ ( .A(_01768_ ), .B1(_01588_ ), .B2(_01644_ ), .ZN(_01769_ ) );
NAND3_X1 _08973_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][19] ), .A3(_01647_ ), .ZN(_01770_ ) );
NAND4_X1 _08974_ ( .A1(_01651_ ), .A2(\u_csr.csr[2][19] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_01771_ ) );
NAND3_X1 _08975_ ( .A1(_01769_ ), .A2(_01770_ ), .A3(_01771_ ), .ZN(_01772_ ) );
NAND3_X1 _08976_ ( .A1(_01439_ ), .A2(_01444_ ), .A3(_01772_ ), .ZN(_01773_ ) );
BUF_X8 _08977_ ( .A(_01472_ ), .Z(_01774_ ) );
NAND4_X1 _08978_ ( .A1(_01774_ ), .A2(_00797_ ), .A3(_00796_ ), .A4(_01715_ ), .ZN(_01775_ ) );
AOI21_X1 _08979_ ( .A(_01767_ ), .B1(_01773_ ), .B2(_01775_ ), .ZN(_01776_ ) );
AOI221_X4 _08980_ ( .A(_01776_ ), .B1(\de_pc [19] ), .B2(_01480_ ), .C1(_01106_ ), .C2(_01109_ ), .ZN(_01777_ ) );
NAND2_X1 _08981_ ( .A1(_01765_ ), .A2(_01485_ ), .ZN(_01778_ ) );
INV_X1 _08982_ ( .A(_01094_ ), .ZN(_01779_ ) );
NOR3_X1 _08983_ ( .A1(_00727_ ), .A2(_00662_ ), .A3(_01779_ ), .ZN(_01780_ ) );
AOI21_X1 _08984_ ( .A(_00662_ ), .B1(_01091_ ), .B2(_00923_ ), .ZN(_01781_ ) );
NOR2_X1 _08985_ ( .A1(_01780_ ), .A2(_01781_ ), .ZN(_01782_ ) );
INV_X1 _08986_ ( .A(_01782_ ), .ZN(_01783_ ) );
NOR2_X1 _08987_ ( .A1(_00721_ ), .A2(_00715_ ), .ZN(_01784_ ) );
INV_X1 _08988_ ( .A(_01784_ ), .ZN(_01785_ ) );
AOI21_X1 _08989_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [19] ), .B2(_01785_ ), .ZN(_01786_ ) );
INV_X1 _08990_ ( .A(_01786_ ), .ZN(_01787_ ) );
AOI221_X1 _08991_ ( .A(_01487_ ), .B1(\de_pc [19] ), .B2(_01492_ ), .C1(_01720_ ), .C2(_01787_ ), .ZN(_01788_ ) );
AOI221_X1 _08992_ ( .A(_00893_ ), .B1(_01766_ ), .B2(_01777_ ), .C1(_01778_ ), .C2(_01788_ ), .ZN(_00133_ ) );
AND3_X1 _08993_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [18] ), .ZN(_01789_ ) );
AOI211_X1 _08994_ ( .A(fanout_net_9 ), .B(_01789_ ), .C1(\ea_addr [18] ), .C2(_01135_ ), .ZN(_01790_ ) );
OR2_X1 _08995_ ( .A1(_01227_ ), .A2(\io_master_rdata [26] ), .ZN(_01791_ ) );
AND3_X1 _08996_ ( .A1(_01212_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ), .A3(_01213_ ), .ZN(_01792_ ) );
INV_X1 _08997_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ), .ZN(_01793_ ) );
OAI21_X1 _08998_ ( .A(_01671_ ), .B1(_01242_ ), .B2(_01793_ ), .ZN(_01794_ ) );
OAI21_X1 _08999_ ( .A(_01526_ ), .B1(_01792_ ), .B2(_01794_ ), .ZN(_01795_ ) );
AND2_X1 _09000_ ( .A1(_01791_ ), .A2(_01795_ ), .ZN(_01796_ ) );
OR2_X1 _09001_ ( .A1(_01796_ ), .A2(_01676_ ), .ZN(_01797_ ) );
OR2_X1 _09002_ ( .A1(_01227_ ), .A2(\io_master_rdata [18] ), .ZN(_01798_ ) );
MUX2_X1 _09003_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ), .B(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ), .S(_01242_ ), .Z(_01799_ ) );
OAI21_X1 _09004_ ( .A(_01526_ ), .B1(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .B2(_01799_ ), .ZN(_01800_ ) );
AOI21_X1 _09005_ ( .A(_01254_ ), .B1(_01798_ ), .B2(_01800_ ), .ZN(_01801_ ) );
NOR4_X1 _09006_ ( .A1(_01801_ ), .A2(\io_master_araddr [1] ), .A3(_01274_ ), .A4(_01275_ ), .ZN(_01802_ ) );
AOI21_X4 _09007_ ( .A(_01273_ ), .B1(_01797_ ), .B2(_01802_ ), .ZN(_01803_ ) );
AOI21_X2 _09008_ ( .A(_01790_ ), .B1(_01803_ ), .B2(fanout_net_9 ), .ZN(\ar_data [18] ) );
NOR2_X1 _09009_ ( .A1(\ar_data [18] ), .A2(_01536_ ), .ZN(_01804_ ) );
BUF_X2 _09010_ ( .A(_01316_ ), .Z(_01805_ ) );
BUF_X4 _09011_ ( .A(_01319_ ), .Z(_01806_ ) );
BUF_X4 _09012_ ( .A(_01758_ ), .Z(_01807_ ) );
AOI22_X1 _09013_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01808_ ) );
BUF_X4 _09014_ ( .A(_01325_ ), .Z(_01809_ ) );
BUF_X4 _09015_ ( .A(_01330_ ), .Z(_01810_ ) );
AOI22_X1 _09016_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01811_ ) );
NAND3_X1 _09017_ ( .A1(_01808_ ), .A2(_01809_ ), .A3(_01811_ ), .ZN(_01812_ ) );
BUF_X4 _09018_ ( .A(_00944_ ), .Z(_01813_ ) );
BUF_X2 _09019_ ( .A(_01813_ ), .Z(_01814_ ) );
OAI211_X1 _09020_ ( .A(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01547_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_01815_ ) );
BUF_X4 _09021_ ( .A(_01694_ ), .Z(_01816_ ) );
INV_X1 _09022_ ( .A(\u_reg.rf[1][18] ), .ZN(_01817_ ) );
AOI21_X1 _09023_ ( .A(_01816_ ), .B1(_01549_ ), .B2(_01817_ ), .ZN(_01818_ ) );
NOR2_X1 _09024_ ( .A1(_01549_ ), .A2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01819_ ) );
OAI211_X1 _09025_ ( .A(_01558_ ), .B(_01815_ ), .C1(_01818_ ), .C2(_01819_ ), .ZN(_01820_ ) );
NAND3_X1 _09026_ ( .A1(_01812_ ), .A2(_01814_ ), .A3(_01820_ ), .ZN(_01821_ ) );
BUF_X2 _09027_ ( .A(_01043_ ), .Z(_01822_ ) );
AOI22_X1 _09028_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01823_ ) );
AOI22_X1 _09029_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01824_ ) );
AOI21_X1 _09030_ ( .A(_01558_ ), .B1(_01823_ ), .B2(_01824_ ), .ZN(_01825_ ) );
AOI22_X1 _09031_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01826_ ) );
AOI22_X1 _09032_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01827_ ) );
AOI21_X1 _09033_ ( .A(_01361_ ), .B1(_01826_ ), .B2(_01827_ ), .ZN(_01828_ ) );
OAI21_X1 _09034_ ( .A(_01822_ ), .B1(_01825_ ), .B2(_01828_ ), .ZN(_01829_ ) );
AOI21_X1 _09035_ ( .A(_01318_ ), .B1(_01821_ ), .B2(_01829_ ), .ZN(_01830_ ) );
OR3_X2 _09036_ ( .A1(_01804_ ), .A2(_01805_ ), .A3(_01830_ ), .ZN(_01831_ ) );
INV_X1 _09037_ ( .A(_00719_ ), .ZN(_01832_ ) );
BUF_X4 _09038_ ( .A(_01832_ ), .Z(_01833_ ) );
NOR2_X1 _09039_ ( .A1(_01831_ ), .A2(_01833_ ), .ZN(_01834_ ) );
AND3_X1 _09040_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][18] ), .A3(_01461_ ), .ZN(_01835_ ) );
AOI21_X1 _09041_ ( .A(_01835_ ), .B1(_01588_ ), .B2(_01644_ ), .ZN(_01836_ ) );
NAND3_X1 _09042_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][18] ), .A3(_01454_ ), .ZN(_01837_ ) );
NAND4_X1 _09043_ ( .A1(_01454_ ), .A2(\u_csr.csr[2][18] ), .A3(_01465_ ), .A4(_01467_ ), .ZN(_01838_ ) );
NAND3_X1 _09044_ ( .A1(_01836_ ), .A2(_01837_ ), .A3(_01838_ ), .ZN(_01839_ ) );
NAND3_X1 _09045_ ( .A1(_01439_ ), .A2(_01444_ ), .A3(_01839_ ), .ZN(_01840_ ) );
NAND4_X1 _09046_ ( .A1(_01774_ ), .A2(_00800_ ), .A3(_00799_ ), .A4(_01443_ ), .ZN(_01841_ ) );
AND2_X1 _09047_ ( .A1(_01840_ ), .A2(_01841_ ), .ZN(_01842_ ) );
BUF_X4 _09048_ ( .A(_01375_ ), .Z(_01843_ ) );
INV_X1 _09049_ ( .A(\de_pc [18] ), .ZN(_01844_ ) );
BUF_X4 _09050_ ( .A(_01478_ ), .Z(_01845_ ) );
OAI22_X1 _09051_ ( .A1(_01842_ ), .A2(_01843_ ), .B1(_01844_ ), .B2(_01845_ ), .ZN(_01846_ ) );
OAI21_X1 _09052_ ( .A(_01070_ ), .B1(_01834_ ), .B2(_01846_ ), .ZN(_01847_ ) );
BUF_X4 _09053_ ( .A(_01483_ ), .Z(_01848_ ) );
BUF_X4 _09054_ ( .A(_01507_ ), .Z(_01849_ ) );
OAI22_X1 _09055_ ( .A1(_01831_ ), .A2(_01848_ ), .B1(_01844_ ), .B2(_01849_ ), .ZN(_01850_ ) );
AOI21_X1 _09056_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [18] ), .B2(_01785_ ), .ZN(_01851_ ) );
INV_X1 _09057_ ( .A(_01851_ ), .ZN(_01852_ ) );
AOI21_X1 _09058_ ( .A(_01850_ ), .B1(_01495_ ), .B2(_01852_ ), .ZN(_01853_ ) );
BUF_X4 _09059_ ( .A(_01570_ ), .Z(_01854_ ) );
OAI21_X1 _09060_ ( .A(_01847_ ), .B1(_01853_ ), .B2(_01854_ ), .ZN(_00134_ ) );
BUF_X4 _09061_ ( .A(_01069_ ), .Z(_01855_ ) );
BUF_X4 _09062_ ( .A(_01313_ ), .Z(_01856_ ) );
AOI22_X1 _09063_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01857_ ) );
BUF_X2 _09064_ ( .A(_01557_ ), .Z(_01858_ ) );
AOI22_X1 _09065_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01859_ ) );
NAND3_X1 _09066_ ( .A1(_01857_ ), .A2(_01858_ ), .A3(_01859_ ), .ZN(_01860_ ) );
AOI22_X1 _09067_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01861_ ) );
AOI22_X1 _09068_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01862_ ) );
NAND3_X1 _09069_ ( .A1(_01861_ ), .A2(_01809_ ), .A3(_01862_ ), .ZN(_01863_ ) );
NAND3_X1 _09070_ ( .A1(_01860_ ), .A2(_01863_ ), .A3(_01822_ ), .ZN(_01864_ ) );
AOI22_X1 _09071_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01865_ ) );
AOI22_X1 _09072_ ( .A1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01866_ ) );
AND3_X1 _09073_ ( .A1(_01865_ ), .A2(_01756_ ), .A3(_01866_ ), .ZN(_01867_ ) );
OR2_X1 _09074_ ( .A1(_01867_ ), .A2(_01366_ ), .ZN(_01868_ ) );
OAI21_X1 _09075_ ( .A(_01338_ ), .B1(_01546_ ), .B2(\u_reg.rf[1][17] ), .ZN(_01869_ ) );
INV_X1 _09076_ ( .A(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01870_ ) );
BUF_X2 _09077_ ( .A(_00933_ ), .Z(_01871_ ) );
BUF_X2 _09078_ ( .A(_00934_ ), .Z(_01872_ ) );
OAI21_X1 _09079_ ( .A(_01870_ ), .B1(_01871_ ), .B2(_01872_ ), .ZN(_01873_ ) );
AOI221_X4 _09080_ ( .A(_01325_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(_01869_ ), .C2(_01873_ ), .ZN(_01874_ ) );
OAI21_X1 _09081_ ( .A(_01864_ ), .B1(_01868_ ), .B2(_01874_ ), .ZN(_01875_ ) );
AOI21_X1 _09082_ ( .A(_01805_ ), .B1(_01856_ ), .B2(_01875_ ), .ZN(_01876_ ) );
AND3_X1 _09083_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [17] ), .ZN(_01877_ ) );
AOI211_X1 _09084_ ( .A(fanout_net_9 ), .B(_01877_ ), .C1(\ea_addr [17] ), .C2(_01135_ ), .ZN(_01878_ ) );
INV_X1 _09085_ ( .A(\u_lsu.u_clint.mtime [17] ), .ZN(_01879_ ) );
NAND4_X1 _09086_ ( .A1(_01239_ ), .A2(_01879_ ), .A3(\io_master_araddr [3] ), .A4(_01266_ ), .ZN(_01880_ ) );
OAI211_X2 _09087_ ( .A(_01238_ ), .B(_01880_ ), .C1(\u_lsu.u_clint.mtime [49] ), .C2(_01733_ ), .ZN(_01881_ ) );
OAI21_X1 _09088_ ( .A(\io_master_rdata [17] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_01882_ ) );
AND3_X1 _09089_ ( .A1(_01881_ ), .A2(_01524_ ), .A3(_01882_ ), .ZN(_01883_ ) );
OR2_X1 _09090_ ( .A1(_01529_ ), .A2(\u_lsu.u_clint.mtime [57] ), .ZN(_01884_ ) );
OAI211_X1 _09091_ ( .A(_01238_ ), .B(_01884_ ), .C1(\u_lsu.u_clint.mtime [25] ), .C2(_01249_ ), .ZN(_01885_ ) );
OAI21_X1 _09092_ ( .A(\io_master_rdata [25] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_01886_ ) );
AND2_X1 _09093_ ( .A1(_01885_ ), .A2(_01886_ ), .ZN(_01887_ ) );
AOI211_X1 _09094_ ( .A(\io_master_araddr [1] ), .B(_01883_ ), .C1(\io_master_araddr [0] ), .C2(_01887_ ), .ZN(_01888_ ) );
AOI21_X2 _09095_ ( .A(_01273_ ), .B1(\io_master_arsize [1] ), .B2(_01888_ ), .ZN(_01889_ ) );
AOI21_X2 _09096_ ( .A(_01878_ ), .B1(_01889_ ), .B2(fanout_net_9 ), .ZN(\ar_data [17] ) );
OAI21_X1 _09097_ ( .A(_01876_ ), .B1(\ar_data [17] ), .B2(_01856_ ), .ZN(_01890_ ) );
NOR2_X1 _09098_ ( .A1(_01890_ ), .A2(_01833_ ), .ZN(_01891_ ) );
NAND4_X1 _09099_ ( .A1(_01455_ ), .A2(\u_csr.csr[2][17] ), .A3(_01653_ ), .A4(_01649_ ), .ZN(_01892_ ) );
NAND3_X1 _09100_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][17] ), .A3(_01455_ ), .ZN(_01893_ ) );
NAND4_X1 _09101_ ( .A1(_01653_ ), .A2(\u_csr.csr[0][17] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_01894_ ) );
NAND4_X1 _09102_ ( .A1(_01646_ ), .A2(_01892_ ), .A3(_01893_ ), .A4(_01894_ ), .ZN(_01895_ ) );
NAND2_X1 _09103_ ( .A1(_01576_ ), .A2(_01895_ ), .ZN(_01896_ ) );
NAND4_X1 _09104_ ( .A1(_01596_ ), .A2(_00802_ ), .A3(_00801_ ), .A4(_01444_ ), .ZN(_01897_ ) );
AND2_X1 _09105_ ( .A1(_01896_ ), .A2(_01897_ ), .ZN(_01898_ ) );
INV_X1 _09106_ ( .A(\de_pc [17] ), .ZN(_01899_ ) );
OAI22_X1 _09107_ ( .A1(_01898_ ), .A2(_01843_ ), .B1(_01899_ ), .B2(_01845_ ), .ZN(_01900_ ) );
OAI21_X1 _09108_ ( .A(_01855_ ), .B1(_01891_ ), .B2(_01900_ ), .ZN(_01901_ ) );
OAI22_X1 _09109_ ( .A1(_01890_ ), .A2(_01848_ ), .B1(_01899_ ), .B2(_01849_ ), .ZN(_01902_ ) );
AOI21_X1 _09110_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [17] ), .B2(_01785_ ), .ZN(_01903_ ) );
INV_X1 _09111_ ( .A(_01903_ ), .ZN(_01904_ ) );
AOI21_X1 _09112_ ( .A(_01902_ ), .B1(_01495_ ), .B2(_01904_ ), .ZN(_01905_ ) );
OAI21_X1 _09113_ ( .A(_01901_ ), .B1(_01905_ ), .B2(_01854_ ), .ZN(_00135_ ) );
AND3_X1 _09114_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [16] ), .ZN(_01906_ ) );
AOI211_X1 _09115_ ( .A(fanout_net_9 ), .B(_01906_ ), .C1(\ea_addr [16] ), .C2(_01136_ ), .ZN(_01907_ ) );
OR2_X1 _09116_ ( .A1(_01527_ ), .A2(\io_master_rdata [24] ), .ZN(_01908_ ) );
BUF_X8 _09117_ ( .A(_01527_ ), .Z(_01909_ ) );
MUX2_X1 _09118_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ), .B(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ), .S(_01529_ ), .Z(_01910_ ) );
OAI21_X1 _09119_ ( .A(_01909_ ), .B1(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .B2(_01910_ ), .ZN(_01911_ ) );
AND2_X1 _09120_ ( .A1(_01908_ ), .A2(_01911_ ), .ZN(_01912_ ) );
OR2_X1 _09121_ ( .A1(_01912_ ), .A2(_01676_ ), .ZN(_01913_ ) );
OR2_X1 _09122_ ( .A1(_01527_ ), .A2(\io_master_rdata [16] ), .ZN(_01914_ ) );
AND3_X1 _09123_ ( .A1(_01669_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ), .A3(_01266_ ), .ZN(_01915_ ) );
INV_X1 _09124_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ), .ZN(_01916_ ) );
OAI21_X1 _09125_ ( .A(_01671_ ), .B1(_01733_ ), .B2(_01916_ ), .ZN(_01917_ ) );
OAI21_X2 _09126_ ( .A(_01909_ ), .B1(_01915_ ), .B2(_01917_ ), .ZN(_01918_ ) );
AOI21_X1 _09127_ ( .A(_01276_ ), .B1(_01914_ ), .B2(_01918_ ), .ZN(_01919_ ) );
NOR4_X1 _09128_ ( .A1(_01919_ ), .A2(\io_master_araddr [1] ), .A3(_01274_ ), .A4(_01275_ ), .ZN(_01920_ ) );
AOI21_X4 _09129_ ( .A(_01273_ ), .B1(_01913_ ), .B2(_01920_ ), .ZN(_01921_ ) );
AOI21_X4 _09130_ ( .A(_01907_ ), .B1(_01921_ ), .B2(fanout_net_9 ), .ZN(\ar_data [16] ) );
NOR2_X2 _09131_ ( .A1(\ar_data [16] ), .A2(_01686_ ), .ZN(_01922_ ) );
AOI22_X1 _09132_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01923_ ) );
AOI22_X1 _09133_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01924_ ) );
NAND3_X1 _09134_ ( .A1(_01923_ ), .A2(_01361_ ), .A3(_01924_ ), .ZN(_01925_ ) );
NAND3_X1 _09135_ ( .A1(_01546_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01338_ ), .ZN(_01926_ ) );
NOR2_X1 _09136_ ( .A1(_01551_ ), .A2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01927_ ) );
BUF_X4 _09137_ ( .A(_01307_ ), .Z(_01928_ ) );
INV_X1 _09138_ ( .A(\u_reg.rf[1][16] ), .ZN(_01929_ ) );
AOI21_X1 _09139_ ( .A(_01694_ ), .B1(_01928_ ), .B2(_01929_ ), .ZN(_01930_ ) );
OAI211_X1 _09140_ ( .A(_01926_ ), .B(_01335_ ), .C1(_01927_ ), .C2(_01930_ ), .ZN(_01931_ ) );
NAND3_X1 _09141_ ( .A1(_01925_ ), .A2(_01334_ ), .A3(_01931_ ), .ZN(_01932_ ) );
AOI22_X1 _09142_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01933_ ) );
AOI22_X1 _09143_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01752_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01934_ ) );
AOI21_X1 _09144_ ( .A(_01557_ ), .B1(_01933_ ), .B2(_01934_ ), .ZN(_01935_ ) );
AOI22_X1 _09145_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01936_ ) );
AOI22_X1 _09146_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01937_ ) );
AOI21_X1 _09147_ ( .A(_01756_ ), .B1(_01936_ ), .B2(_01937_ ), .ZN(_01938_ ) );
OAI21_X1 _09148_ ( .A(_01366_ ), .B1(_01935_ ), .B2(_01938_ ), .ZN(_01939_ ) );
AOI21_X1 _09149_ ( .A(_01688_ ), .B1(_01932_ ), .B2(_01939_ ), .ZN(_01940_ ) );
NOR3_X2 _09150_ ( .A1(_01922_ ), .A2(_01317_ ), .A3(_01940_ ), .ZN(_01941_ ) );
NAND2_X1 _09151_ ( .A1(_01941_ ), .A2(_01371_ ), .ZN(_01942_ ) );
AND3_X1 _09152_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][16] ), .A3(_01647_ ), .ZN(_01943_ ) );
AND3_X1 _09153_ ( .A1(_01457_ ), .A2(\u_csr.csr[0][16] ), .A3(_01460_ ), .ZN(_01944_ ) );
AOI21_X1 _09154_ ( .A(_01944_ ), .B1(_01583_ ), .B2(_01587_ ), .ZN(_01945_ ) );
NAND4_X1 _09155_ ( .A1(_01582_ ), .A2(\u_csr.csr[2][16] ), .A3(_00754_ ), .A4(_01591_ ), .ZN(_01946_ ) );
NAND2_X1 _09156_ ( .A1(_01945_ ), .A2(_01946_ ), .ZN(_01947_ ) );
OAI21_X1 _09157_ ( .A(_01575_ ), .B1(_01943_ ), .B2(_01947_ ), .ZN(_01948_ ) );
NAND4_X1 _09158_ ( .A1(_01774_ ), .A2(_00804_ ), .A3(_00803_ ), .A4(_01715_ ), .ZN(_01949_ ) );
AOI21_X1 _09159_ ( .A(_01767_ ), .B1(_01948_ ), .B2(_01949_ ), .ZN(_01950_ ) );
AOI221_X4 _09160_ ( .A(_01950_ ), .B1(\de_pc [16] ), .B2(_01480_ ), .C1(_01106_ ), .C2(_01109_ ), .ZN(_01951_ ) );
NAND2_X1 _09161_ ( .A1(_01941_ ), .A2(_01485_ ), .ZN(_01952_ ) );
AOI21_X1 _09162_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [16] ), .B2(_01785_ ), .ZN(_01953_ ) );
INV_X1 _09163_ ( .A(_01953_ ), .ZN(_01954_ ) );
AOI221_X1 _09164_ ( .A(_01487_ ), .B1(\de_pc [16] ), .B2(_01492_ ), .C1(_01720_ ), .C2(_01954_ ), .ZN(_01955_ ) );
AOI221_X1 _09165_ ( .A(_00893_ ), .B1(_01942_ ), .B2(_01951_ ), .C1(_01952_ ), .C2(_01955_ ), .ZN(_00136_ ) );
AND3_X1 _09166_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [15] ), .ZN(_01956_ ) );
AOI211_X1 _09167_ ( .A(fanout_net_9 ), .B(_01956_ ), .C1(\ea_addr [15] ), .C2(_01135_ ), .ZN(_01957_ ) );
INV_X1 _09168_ ( .A(_01274_ ), .ZN(_01958_ ) );
AOI21_X2 _09169_ ( .A(_01604_ ), .B1(_01958_ ), .B2(_01269_ ), .ZN(_01959_ ) );
AOI21_X2 _09170_ ( .A(_01957_ ), .B1(_01959_ ), .B2(fanout_net_9 ), .ZN(\ar_data [15] ) );
NOR2_X1 _09171_ ( .A1(\ar_data [15] ), .A2(_01536_ ), .ZN(_01960_ ) );
AOI22_X1 _09172_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01961_ ) );
AOI22_X1 _09173_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01962_ ) );
NAND3_X1 _09174_ ( .A1(_01961_ ), .A2(_01809_ ), .A3(_01962_ ), .ZN(_01963_ ) );
BUF_X4 _09175_ ( .A(_01545_ ), .Z(_01964_ ) );
BUF_X4 _09176_ ( .A(_01337_ ), .Z(_01965_ ) );
NAND3_X1 _09177_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01965_ ), .ZN(_01966_ ) );
NOR2_X1 _09178_ ( .A1(_01549_ ), .A2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01967_ ) );
INV_X1 _09179_ ( .A(\u_reg.rf[1][15] ), .ZN(_01968_ ) );
AOI21_X1 _09180_ ( .A(_01343_ ), .B1(_01549_ ), .B2(_01968_ ), .ZN(_01969_ ) );
OAI211_X1 _09181_ ( .A(_01966_ ), .B(_01558_ ), .C1(_01967_ ), .C2(_01969_ ), .ZN(_01970_ ) );
NAND3_X1 _09182_ ( .A1(_01963_ ), .A2(_01814_ ), .A3(_01970_ ), .ZN(_01971_ ) );
AOI22_X1 _09183_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01972_ ) );
AOI22_X1 _09184_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01973_ ) );
AOI21_X1 _09185_ ( .A(_01558_ ), .B1(_01972_ ), .B2(_01973_ ), .ZN(_01974_ ) );
AOI22_X1 _09186_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01975_ ) );
AOI22_X1 _09187_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01976_ ) );
AOI21_X1 _09188_ ( .A(_01361_ ), .B1(_01975_ ), .B2(_01976_ ), .ZN(_01977_ ) );
OAI21_X1 _09189_ ( .A(_01822_ ), .B1(_01974_ ), .B2(_01977_ ), .ZN(_01978_ ) );
AOI21_X1 _09190_ ( .A(_01318_ ), .B1(_01971_ ), .B2(_01978_ ), .ZN(_01979_ ) );
OR3_X2 _09191_ ( .A1(_01960_ ), .A2(_01805_ ), .A3(_01979_ ), .ZN(_01980_ ) );
NOR2_X1 _09192_ ( .A1(_01980_ ), .A2(_01833_ ), .ZN(_01981_ ) );
NAND3_X1 _09193_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][15] ), .A3(_01455_ ), .ZN(_01982_ ) );
NAND3_X1 _09194_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][15] ), .A3(_01461_ ), .ZN(_01983_ ) );
NAND4_X1 _09195_ ( .A1(_01454_ ), .A2(\u_csr.csr[2][15] ), .A3(_01465_ ), .A4(_01467_ ), .ZN(_01984_ ) );
NAND3_X1 _09196_ ( .A1(_01982_ ), .A2(_01983_ ), .A3(_01984_ ), .ZN(_01985_ ) );
NAND3_X1 _09197_ ( .A1(_01439_ ), .A2(_01715_ ), .A3(_01985_ ), .ZN(_01986_ ) );
NAND4_X1 _09198_ ( .A1(_01472_ ), .A2(_00807_ ), .A3(_00805_ ), .A4(_01443_ ), .ZN(_01987_ ) );
AND2_X1 _09199_ ( .A1(_01986_ ), .A2(_01987_ ), .ZN(_01988_ ) );
INV_X1 _09200_ ( .A(\de_pc [15] ), .ZN(_01989_ ) );
OAI22_X1 _09201_ ( .A1(_01988_ ), .A2(_01843_ ), .B1(_01989_ ), .B2(_01845_ ), .ZN(_01990_ ) );
OAI21_X1 _09202_ ( .A(_01855_ ), .B1(_01981_ ), .B2(_01990_ ), .ZN(_01991_ ) );
OAI22_X1 _09203_ ( .A1(_01980_ ), .A2(_01848_ ), .B1(_01989_ ), .B2(_01849_ ), .ZN(_01992_ ) );
AOI21_X1 _09204_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [15] ), .B2(_01785_ ), .ZN(_01993_ ) );
INV_X1 _09205_ ( .A(_01993_ ), .ZN(_01994_ ) );
AOI21_X1 _09206_ ( .A(_01992_ ), .B1(_01495_ ), .B2(_01994_ ), .ZN(_01995_ ) );
OAI21_X1 _09207_ ( .A(_01991_ ), .B1(_01995_ ), .B2(_01854_ ), .ZN(_00137_ ) );
AND3_X1 _09208_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [14] ), .ZN(_01996_ ) );
AOI211_X1 _09209_ ( .A(fanout_net_9 ), .B(_01996_ ), .C1(\ea_addr [14] ), .C2(_01136_ ), .ZN(_01997_ ) );
OR2_X1 _09210_ ( .A1(_01527_ ), .A2(\io_master_rdata [22] ), .ZN(_01998_ ) );
AND3_X1 _09211_ ( .A1(_01669_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_39_A_$_ANDNOT__Y_B ), .A3(_01266_ ), .ZN(_01999_ ) );
INV_X1 _09212_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_8_A_$_ANDNOT__Y_B ), .ZN(_02000_ ) );
OAI21_X1 _09213_ ( .A(_01671_ ), .B1(_01733_ ), .B2(_02000_ ), .ZN(_02001_ ) );
OAI21_X1 _09214_ ( .A(_01527_ ), .B1(_01999_ ), .B2(_02001_ ), .ZN(_02002_ ) );
AND3_X1 _09215_ ( .A1(_01998_ ), .A2(_01143_ ), .A3(_02002_ ), .ZN(_02003_ ) );
BUF_X2 _09216_ ( .A(_01246_ ), .Z(_02004_ ) );
AOI21_X1 _09217_ ( .A(_02003_ ), .B1(_02004_ ), .B2(_01532_ ), .ZN(_02005_ ) );
MUX2_X1 _09218_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ), .B(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ), .S(_01733_ ), .Z(_02006_ ) );
OAI21_X1 _09219_ ( .A(_01909_ ), .B1(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .B2(_02006_ ), .ZN(_02007_ ) );
OAI21_X1 _09220_ ( .A(_02007_ ), .B1(\io_master_rdata [14] ), .B2(_01909_ ), .ZN(_02008_ ) );
OAI21_X1 _09221_ ( .A(_02005_ ), .B1(_01277_ ), .B2(_02008_ ), .ZN(_02009_ ) );
AOI21_X2 _09222_ ( .A(_01604_ ), .B1(_01958_ ), .B2(_02009_ ), .ZN(_02010_ ) );
AOI21_X2 _09223_ ( .A(_01997_ ), .B1(_02010_ ), .B2(fanout_net_9 ), .ZN(\ar_data [14] ) );
OR2_X1 _09224_ ( .A1(\ar_data [14] ), .A2(_01536_ ), .ZN(_02011_ ) );
BUF_X4 _09225_ ( .A(_01749_ ), .Z(_02012_ ) );
BUF_X4 _09226_ ( .A(_01750_ ), .Z(_02013_ ) );
AOI22_X1 _09227_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_02012_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02014_ ) );
BUF_X2 _09228_ ( .A(_01325_ ), .Z(_02015_ ) );
BUF_X4 _09229_ ( .A(_01752_ ), .Z(_02016_ ) );
BUF_X4 _09230_ ( .A(_01760_ ), .Z(_02017_ ) );
AOI22_X1 _09231_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02018_ ) );
NAND3_X1 _09232_ ( .A1(_02014_ ), .A2(_02015_ ), .A3(_02018_ ), .ZN(_02019_ ) );
NAND3_X1 _09233_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01965_ ), .ZN(_02020_ ) );
BUF_X4 _09234_ ( .A(_01928_ ), .Z(_02021_ ) );
NOR2_X1 _09235_ ( .A1(_02021_ ), .A2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02022_ ) );
INV_X1 _09236_ ( .A(\u_reg.rf[1][14] ), .ZN(_02023_ ) );
AOI21_X1 _09237_ ( .A(_01816_ ), .B1(_01549_ ), .B2(_02023_ ), .ZN(_02024_ ) );
OAI211_X1 _09238_ ( .A(_02020_ ), .B(_01858_ ), .C1(_02022_ ), .C2(_02024_ ), .ZN(_02025_ ) );
AND3_X1 _09239_ ( .A1(_02019_ ), .A2(_01814_ ), .A3(_02025_ ), .ZN(_02026_ ) );
AOI22_X1 _09240_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02027_ ) );
AOI22_X1 _09241_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02028_ ) );
NAND3_X1 _09242_ ( .A1(_02027_ ), .A2(_01858_ ), .A3(_02028_ ), .ZN(_02029_ ) );
AOI22_X1 _09243_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02030_ ) );
AOI22_X1 _09244_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02031_ ) );
NAND3_X1 _09245_ ( .A1(_02030_ ), .A2(_02015_ ), .A3(_02031_ ), .ZN(_02032_ ) );
AND3_X1 _09246_ ( .A1(_02029_ ), .A2(_02032_ ), .A3(_01822_ ), .ZN(_02033_ ) );
OAI21_X1 _09247_ ( .A(_01856_ ), .B1(_02026_ ), .B2(_02033_ ), .ZN(_02034_ ) );
NAND3_X1 _09248_ ( .A1(_02011_ ), .A2(_01535_ ), .A3(_02034_ ), .ZN(_02035_ ) );
NOR2_X1 _09249_ ( .A1(_02035_ ), .A2(_01833_ ), .ZN(_02036_ ) );
AND3_X1 _09250_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][14] ), .A3(_01455_ ), .ZN(_02037_ ) );
AND3_X1 _09251_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][14] ), .A3(_01461_ ), .ZN(_02038_ ) );
AOI21_X1 _09252_ ( .A(_02038_ ), .B1(_01583_ ), .B2(_01588_ ), .ZN(_02039_ ) );
NAND4_X1 _09253_ ( .A1(_01583_ ), .A2(\u_csr.csr[2][14] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_02040_ ) );
NAND2_X1 _09254_ ( .A1(_02039_ ), .A2(_02040_ ), .ZN(_02041_ ) );
OAI21_X1 _09255_ ( .A(_01576_ ), .B1(_02037_ ), .B2(_02041_ ), .ZN(_02042_ ) );
NAND4_X1 _09256_ ( .A1(_01596_ ), .A2(_00809_ ), .A3(_00808_ ), .A4(_01444_ ), .ZN(_02043_ ) );
AND2_X1 _09257_ ( .A1(_02042_ ), .A2(_02043_ ), .ZN(_02044_ ) );
INV_X1 _09258_ ( .A(\de_pc [14] ), .ZN(_02045_ ) );
OAI22_X1 _09259_ ( .A1(_02044_ ), .A2(_01843_ ), .B1(_02045_ ), .B2(_01845_ ), .ZN(_02046_ ) );
OAI21_X1 _09260_ ( .A(_01855_ ), .B1(_02036_ ), .B2(_02046_ ), .ZN(_02047_ ) );
OAI22_X1 _09261_ ( .A1(_02035_ ), .A2(_01848_ ), .B1(_02045_ ), .B2(_01849_ ), .ZN(_02048_ ) );
AOI21_X1 _09262_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [14] ), .B2(_01785_ ), .ZN(_02049_ ) );
INV_X1 _09263_ ( .A(_02049_ ), .ZN(_02050_ ) );
AOI21_X1 _09264_ ( .A(_02048_ ), .B1(_01495_ ), .B2(_02050_ ), .ZN(_02051_ ) );
OAI21_X1 _09265_ ( .A(_02047_ ), .B1(_02051_ ), .B2(_01854_ ), .ZN(_00138_ ) );
AND3_X1 _09266_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [13] ), .ZN(_02052_ ) );
AOI211_X1 _09267_ ( .A(fanout_net_9 ), .B(_02052_ ), .C1(\ea_addr [13] ), .C2(_01136_ ), .ZN(_02053_ ) );
INV_X1 _09268_ ( .A(_01669_ ), .ZN(_02054_ ) );
NOR3_X1 _09269_ ( .A1(_02054_ ), .A2(\u_lsu.u_clint.mtime [13] ), .A3(_01254_ ), .ZN(_02055_ ) );
INV_X1 _09270_ ( .A(\u_lsu.u_clint.mtime [45] ), .ZN(_02056_ ) );
AOI211_X2 _09271_ ( .A(_02055_ ), .B(_01229_ ), .C1(_02056_ ), .C2(_01249_ ), .ZN(_02057_ ) );
INV_X4 _09272_ ( .A(_01526_ ), .ZN(io_master_rready ) );
AND2_X1 _09273_ ( .A1(io_master_rready ), .A2(\io_master_rdata [13] ), .ZN(_02058_ ) );
NOR3_X1 _09274_ ( .A1(_02057_ ), .A2(_01254_ ), .A3(_02058_ ), .ZN(_02059_ ) );
AOI21_X1 _09275_ ( .A(_01144_ ), .B1(_01606_ ), .B2(_01609_ ), .ZN(_02060_ ) );
AOI21_X1 _09276_ ( .A(_02060_ ), .B1(_02004_ ), .B2(_01614_ ), .ZN(_02061_ ) );
AOI211_X1 _09277_ ( .A(_01274_ ), .B(_02059_ ), .C1(_01276_ ), .C2(_02061_ ), .ZN(_02062_ ) );
NOR2_X2 _09278_ ( .A1(_01604_ ), .A2(_02062_ ), .ZN(_02063_ ) );
AOI21_X2 _09279_ ( .A(_02053_ ), .B1(_02063_ ), .B2(fanout_net_9 ), .ZN(\ar_data [13] ) );
OR2_X1 _09280_ ( .A1(\ar_data [13] ), .A2(_01536_ ), .ZN(_02064_ ) );
AOI22_X1 _09281_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_02012_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02065_ ) );
AOI22_X1 _09282_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02066_ ) );
NAND3_X1 _09283_ ( .A1(_02065_ ), .A2(_02015_ ), .A3(_02066_ ), .ZN(_02067_ ) );
NAND3_X1 _09284_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01965_ ), .ZN(_02068_ ) );
NOR2_X1 _09285_ ( .A1(_02021_ ), .A2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02069_ ) );
INV_X1 _09286_ ( .A(\u_reg.rf[1][13] ), .ZN(_02070_ ) );
AOI21_X1 _09287_ ( .A(_01816_ ), .B1(_01549_ ), .B2(_02070_ ), .ZN(_02071_ ) );
OAI211_X1 _09288_ ( .A(_02068_ ), .B(_01858_ ), .C1(_02069_ ), .C2(_02071_ ), .ZN(_02072_ ) );
AND3_X1 _09289_ ( .A1(_02067_ ), .A2(_01814_ ), .A3(_02072_ ), .ZN(_02073_ ) );
AOI22_X1 _09290_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02074_ ) );
AOI22_X1 _09291_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02075_ ) );
NAND3_X1 _09292_ ( .A1(_02074_ ), .A2(_01858_ ), .A3(_02075_ ), .ZN(_02076_ ) );
AOI22_X1 _09293_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02077_ ) );
AOI22_X1 _09294_ ( .A1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02078_ ) );
NAND3_X1 _09295_ ( .A1(_02077_ ), .A2(_02015_ ), .A3(_02078_ ), .ZN(_02079_ ) );
AND3_X1 _09296_ ( .A1(_02076_ ), .A2(_02079_ ), .A3(_01822_ ), .ZN(_02080_ ) );
OAI21_X1 _09297_ ( .A(_01856_ ), .B1(_02073_ ), .B2(_02080_ ), .ZN(_02081_ ) );
NAND3_X1 _09298_ ( .A1(_02064_ ), .A2(_01535_ ), .A3(_02081_ ), .ZN(_02082_ ) );
NOR2_X1 _09299_ ( .A1(_02082_ ), .A2(_01833_ ), .ZN(_02083_ ) );
AND3_X1 _09300_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][13] ), .A3(_01461_ ), .ZN(_02084_ ) );
AOI21_X1 _09301_ ( .A(_02084_ ), .B1(_01583_ ), .B2(_01587_ ), .ZN(_02085_ ) );
NAND3_X1 _09302_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][13] ), .A3(_01454_ ), .ZN(_02086_ ) );
NAND4_X1 _09303_ ( .A1(_01454_ ), .A2(\u_csr.csr[2][13] ), .A3(_01465_ ), .A4(_01467_ ), .ZN(_02087_ ) );
NAND3_X1 _09304_ ( .A1(_02085_ ), .A2(_02086_ ), .A3(_02087_ ), .ZN(_02088_ ) );
NAND3_X1 _09305_ ( .A1(_01439_ ), .A2(_01715_ ), .A3(_02088_ ), .ZN(_02089_ ) );
NAND4_X1 _09306_ ( .A1(_01472_ ), .A2(_00811_ ), .A3(_00810_ ), .A4(_01443_ ), .ZN(_02090_ ) );
AND2_X1 _09307_ ( .A1(_02089_ ), .A2(_02090_ ), .ZN(_02091_ ) );
INV_X1 _09308_ ( .A(\de_pc [13] ), .ZN(_02092_ ) );
OAI22_X1 _09309_ ( .A1(_02091_ ), .A2(_01843_ ), .B1(_02092_ ), .B2(_01845_ ), .ZN(_02093_ ) );
OAI21_X1 _09310_ ( .A(_01855_ ), .B1(_02083_ ), .B2(_02093_ ), .ZN(_02094_ ) );
OAI22_X1 _09311_ ( .A1(_02082_ ), .A2(_01848_ ), .B1(_02092_ ), .B2(_01849_ ), .ZN(_02095_ ) );
AOI21_X1 _09312_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [13] ), .B2(_01785_ ), .ZN(_02096_ ) );
INV_X1 _09313_ ( .A(_02096_ ), .ZN(_02097_ ) );
AOI21_X1 _09314_ ( .A(_02095_ ), .B1(_01495_ ), .B2(_02097_ ), .ZN(_02098_ ) );
OAI21_X1 _09315_ ( .A(_02094_ ), .B1(_02098_ ), .B2(_01854_ ), .ZN(_00139_ ) );
AND3_X1 _09316_ ( .A1(_01678_ ), .A2(_01143_ ), .A3(_01682_ ), .ZN(_02099_ ) );
AOI21_X1 _09317_ ( .A(_02099_ ), .B1(_02004_ ), .B2(_01675_ ), .ZN(_02100_ ) );
AND3_X1 _09318_ ( .A1(_01669_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ), .A3(_01266_ ), .ZN(_02101_ ) );
INV_X1 _09319_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_18_A_$_ANDNOT__Y_B ), .ZN(_02102_ ) );
OAI21_X1 _09320_ ( .A(_01671_ ), .B1(_01733_ ), .B2(_02102_ ), .ZN(_02103_ ) );
OAI21_X1 _09321_ ( .A(_01909_ ), .B1(_02101_ ), .B2(_02103_ ), .ZN(_02104_ ) );
OAI21_X1 _09322_ ( .A(_02104_ ), .B1(\io_master_rdata [12] ), .B2(_01909_ ), .ZN(_02105_ ) );
OAI21_X1 _09323_ ( .A(_02100_ ), .B1(_01276_ ), .B2(_02105_ ), .ZN(_02106_ ) );
AOI21_X1 _09324_ ( .A(_01263_ ), .B1(_01958_ ), .B2(_02106_ ), .ZN(_02107_ ) );
NAND2_X1 _09325_ ( .A1(_02107_ ), .A2(fanout_net_9 ), .ZN(_02108_ ) );
MUX2_X1 _09326_ ( .A(\u_exu.ecsr [12] ), .B(\ea_addr [12] ), .S(_01134_ ), .Z(_02109_ ) );
OR2_X1 _09327_ ( .A1(_02109_ ), .A2(fanout_net_9 ), .ZN(_02110_ ) );
AOI21_X1 _09328_ ( .A(_01686_ ), .B1(_02108_ ), .B2(_02110_ ), .ZN(_02111_ ) );
AOI22_X1 _09329_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01017_ ), .B1(_01321_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02112_ ) );
AOI22_X1 _09330_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01327_ ), .B1(_01329_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02113_ ) );
AND3_X1 _09331_ ( .A1(_02112_ ), .A2(_01324_ ), .A3(_02113_ ), .ZN(_02114_ ) );
OAI21_X1 _09332_ ( .A(_01336_ ), .B1(_01292_ ), .B2(\u_reg.rf[1][12] ), .ZN(_02115_ ) );
OR2_X1 _09333_ ( .A1(_01307_ ), .A2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02116_ ) );
AOI221_X4 _09334_ ( .A(_01324_ ), .B1(_01329_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(_02115_ ), .C2(_02116_ ), .ZN(_02117_ ) );
OR3_X1 _09335_ ( .A1(_02114_ ), .A2(_01043_ ), .A3(_02117_ ), .ZN(_02118_ ) );
AOI22_X1 _09336_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02119_ ) );
AOI22_X1 _09337_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02120_ ) );
NAND3_X1 _09338_ ( .A1(_02119_ ), .A2(_01354_ ), .A3(_02120_ ), .ZN(_02121_ ) );
AOI22_X1 _09339_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02122_ ) );
AOI22_X1 _09340_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02123_ ) );
NAND3_X1 _09341_ ( .A1(_02122_ ), .A2(_01633_ ), .A3(_02123_ ), .ZN(_02124_ ) );
NAND3_X1 _09342_ ( .A1(_02121_ ), .A2(_02124_ ), .A3(_01705_ ), .ZN(_02125_ ) );
AOI21_X1 _09343_ ( .A(_01688_ ), .B1(_02118_ ), .B2(_02125_ ), .ZN(_02126_ ) );
NOR3_X1 _09344_ ( .A1(_02111_ ), .A2(_01317_ ), .A3(_02126_ ), .ZN(_02127_ ) );
NAND2_X1 _09345_ ( .A1(_02127_ ), .A2(_01371_ ), .ZN(_02128_ ) );
AND2_X1 _09346_ ( .A1(_01472_ ), .A2(_01442_ ), .ZN(_02129_ ) );
OR2_X1 _09347_ ( .A1(\ea_addr [12] ), .A2(ea_err ), .ZN(_02130_ ) );
OAI211_X1 _09348_ ( .A(_02129_ ), .B(_02130_ ), .C1(_00788_ ), .C2(\ea_pc [12] ), .ZN(_02131_ ) );
NAND4_X1 _09349_ ( .A1(_01651_ ), .A2(\u_csr.csr[2][12] ), .A3(_01465_ ), .A4(_01467_ ), .ZN(_02132_ ) );
NAND3_X1 _09350_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][12] ), .A3(_01454_ ), .ZN(_02133_ ) );
NAND4_X1 _09351_ ( .A1(_01648_ ), .A2(\u_csr.csr[0][12] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_02134_ ) );
NAND4_X1 _09352_ ( .A1(_01646_ ), .A2(_02132_ ), .A3(_02133_ ), .A4(_02134_ ), .ZN(_02135_ ) );
NAND2_X1 _09353_ ( .A1(_01575_ ), .A2(_02135_ ), .ZN(_02136_ ) );
AOI21_X1 _09354_ ( .A(_01767_ ), .B1(_02131_ ), .B2(_02136_ ), .ZN(_02137_ ) );
AOI221_X1 _09355_ ( .A(_02137_ ), .B1(\de_pc [12] ), .B2(_01480_ ), .C1(_01106_ ), .C2(_01109_ ), .ZN(_02138_ ) );
NAND2_X1 _09356_ ( .A1(_02127_ ), .A2(_01485_ ), .ZN(_02139_ ) );
AOI21_X1 _09357_ ( .A(_01783_ ), .B1(\u_idu.imm_auipc_lui [12] ), .B2(_01785_ ), .ZN(_02140_ ) );
INV_X1 _09358_ ( .A(_02140_ ), .ZN(_02141_ ) );
AOI221_X1 _09359_ ( .A(_01487_ ), .B1(\de_pc [12] ), .B2(_01491_ ), .C1(_01720_ ), .C2(_02141_ ), .ZN(_02142_ ) );
AOI221_X1 _09360_ ( .A(_00893_ ), .B1(_02128_ ), .B2(_02138_ ), .C1(_02139_ ), .C2(_02142_ ), .ZN(_00140_ ) );
AND3_X1 _09361_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [29] ), .ZN(_02143_ ) );
AOI211_X1 _09362_ ( .A(fanout_net_9 ), .B(_02143_ ), .C1(\ea_addr [29] ), .C2(_01521_ ), .ZN(_02144_ ) );
AOI21_X2 _09363_ ( .A(_01523_ ), .B1(_01525_ ), .B2(_01614_ ), .ZN(_02145_ ) );
AOI21_X2 _09364_ ( .A(_02144_ ), .B1(_02145_ ), .B2(fanout_net_10 ), .ZN(\ar_data [29] ) );
NOR2_X2 _09365_ ( .A1(\ar_data [29] ), .A2(_01686_ ), .ZN(_02146_ ) );
AOI22_X1 _09366_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02147_ ) );
AOI22_X1 _09367_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02148_ ) );
NAND3_X1 _09368_ ( .A1(_02147_ ), .A2(_01361_ ), .A3(_02148_ ), .ZN(_02149_ ) );
NAND3_X1 _09369_ ( .A1(_01546_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01338_ ), .ZN(_02150_ ) );
NOR2_X1 _09370_ ( .A1(_01551_ ), .A2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02151_ ) );
INV_X1 _09371_ ( .A(\u_reg.rf[1][29] ), .ZN(_02152_ ) );
AOI21_X1 _09372_ ( .A(_01694_ ), .B1(_01928_ ), .B2(_02152_ ), .ZN(_02153_ ) );
OAI211_X1 _09373_ ( .A(_02150_ ), .B(_01557_ ), .C1(_02151_ ), .C2(_02153_ ), .ZN(_02154_ ) );
NAND3_X1 _09374_ ( .A1(_02149_ ), .A2(_01813_ ), .A3(_02154_ ), .ZN(_02155_ ) );
AOI22_X1 _09375_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02156_ ) );
AOI22_X1 _09376_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02157_ ) );
NAND3_X1 _09377_ ( .A1(_02156_ ), .A2(_01354_ ), .A3(_02157_ ), .ZN(_02158_ ) );
AOI22_X1 _09378_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02159_ ) );
AOI22_X1 _09379_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02160_ ) );
NAND3_X1 _09380_ ( .A1(_02159_ ), .A2(_01633_ ), .A3(_02160_ ), .ZN(_02161_ ) );
NAND3_X1 _09381_ ( .A1(_02158_ ), .A2(_02161_ ), .A3(_01705_ ), .ZN(_02162_ ) );
AOI21_X1 _09382_ ( .A(_01688_ ), .B1(_02155_ ), .B2(_02162_ ), .ZN(_02163_ ) );
NOR3_X2 _09383_ ( .A1(_02146_ ), .A2(_01317_ ), .A3(_02163_ ), .ZN(_02164_ ) );
NAND2_X1 _09384_ ( .A1(_02164_ ), .A2(_01370_ ), .ZN(_02165_ ) );
AND3_X1 _09385_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][29] ), .A3(_01461_ ), .ZN(_02166_ ) );
AOI21_X1 _09386_ ( .A(_02166_ ), .B1(_01583_ ), .B2(_01587_ ), .ZN(_02167_ ) );
NAND3_X1 _09387_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][29] ), .A3(_01647_ ), .ZN(_02168_ ) );
NAND4_X1 _09388_ ( .A1(_01651_ ), .A2(\u_csr.csr[2][29] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_02169_ ) );
NAND3_X1 _09389_ ( .A1(_02167_ ), .A2(_02168_ ), .A3(_02169_ ), .ZN(_02170_ ) );
NAND3_X1 _09390_ ( .A1(_01439_ ), .A2(_01444_ ), .A3(_02170_ ), .ZN(_02171_ ) );
NAND4_X1 _09391_ ( .A1(_01774_ ), .A2(_00815_ ), .A3(_00814_ ), .A4(_01715_ ), .ZN(_02172_ ) );
AOI21_X1 _09392_ ( .A(_01767_ ), .B1(_02171_ ), .B2(_02172_ ), .ZN(_02173_ ) );
AOI221_X4 _09393_ ( .A(_02173_ ), .B1(\de_pc [29] ), .B2(_01480_ ), .C1(_01106_ ), .C2(_01108_ ), .ZN(_02174_ ) );
NAND2_X1 _09394_ ( .A1(_02164_ ), .A2(_01484_ ), .ZN(_02175_ ) );
NAND3_X1 _09395_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [29] ), .A3(_01512_ ), .ZN(_02176_ ) );
AND3_X1 _09396_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_02176_ ), .ZN(_02177_ ) );
NOR2_X1 _09397_ ( .A1(_01509_ ), .A2(_02177_ ), .ZN(_02178_ ) );
AOI211_X1 _09398_ ( .A(_02178_ ), .B(_01057_ ), .C1(\de_pc [29] ), .C2(_01492_ ), .ZN(_02179_ ) );
AOI221_X1 _09399_ ( .A(_00893_ ), .B1(_02165_ ), .B2(_02174_ ), .C1(_02175_ ), .C2(_02179_ ), .ZN(_00141_ ) );
AND3_X1 _09400_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [11] ), .ZN(_02180_ ) );
AOI211_X1 _09401_ ( .A(fanout_net_10 ), .B(_02180_ ), .C1(\ea_addr [11] ), .C2(_01521_ ), .ZN(_02181_ ) );
AOI21_X1 _09402_ ( .A(_01144_ ), .B1(_01728_ ), .B2(_01729_ ), .ZN(_02182_ ) );
AOI21_X1 _09403_ ( .A(_02182_ ), .B1(_02004_ ), .B2(_01736_ ), .ZN(_02183_ ) );
AOI21_X1 _09404_ ( .A(\u_lsu.u_clint.mtime [43] ), .B1(_01212_ ), .B2(_01213_ ), .ZN(_02184_ ) );
INV_X1 _09405_ ( .A(\u_lsu.u_clint.mtime [11] ), .ZN(_02185_ ) );
AOI211_X2 _09406_ ( .A(_02184_ ), .B(_01229_ ), .C1(_02185_ ), .C2(_01242_ ), .ZN(_02186_ ) );
AOI21_X2 _09407_ ( .A(_02186_ ), .B1(\io_master_rdata [11] ), .B2(io_master_rready ), .ZN(_02187_ ) );
OAI21_X1 _09408_ ( .A(_02183_ ), .B1(_02187_ ), .B2(_01277_ ), .ZN(_02188_ ) );
AOI21_X2 _09409_ ( .A(_01604_ ), .B1(_01958_ ), .B2(_02188_ ), .ZN(_02189_ ) );
AOI21_X2 _09410_ ( .A(_02181_ ), .B1(_02189_ ), .B2(fanout_net_10 ), .ZN(\ar_data [11] ) );
NOR2_X1 _09411_ ( .A1(\ar_data [11] ), .A2(_01313_ ), .ZN(_02190_ ) );
AOI22_X1 _09412_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02191_ ) );
AOI22_X1 _09413_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02192_ ) );
NAND3_X1 _09414_ ( .A1(_02191_ ), .A2(_01809_ ), .A3(_02192_ ), .ZN(_02193_ ) );
NAND3_X1 _09415_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01965_ ), .ZN(_02194_ ) );
NOR2_X1 _09416_ ( .A1(_01549_ ), .A2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02195_ ) );
INV_X1 _09417_ ( .A(\u_reg.rf[1][11] ), .ZN(_02196_ ) );
AOI21_X1 _09418_ ( .A(_01343_ ), .B1(_01549_ ), .B2(_02196_ ), .ZN(_02197_ ) );
OAI211_X1 _09419_ ( .A(_02194_ ), .B(_01558_ ), .C1(_02195_ ), .C2(_02197_ ), .ZN(_02198_ ) );
NAND3_X1 _09420_ ( .A1(_02193_ ), .A2(_01814_ ), .A3(_02198_ ), .ZN(_02199_ ) );
AOI22_X1 _09421_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02200_ ) );
AOI22_X1 _09422_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02201_ ) );
AOI21_X1 _09423_ ( .A(_01558_ ), .B1(_02200_ ), .B2(_02201_ ), .ZN(_02202_ ) );
AOI22_X1 _09424_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02203_ ) );
AOI22_X1 _09425_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02204_ ) );
AOI21_X1 _09426_ ( .A(_01361_ ), .B1(_02203_ ), .B2(_02204_ ), .ZN(_02205_ ) );
OAI21_X1 _09427_ ( .A(_01822_ ), .B1(_02202_ ), .B2(_02205_ ), .ZN(_02206_ ) );
AOI21_X1 _09428_ ( .A(_01318_ ), .B1(_02199_ ), .B2(_02206_ ), .ZN(_02207_ ) );
OR3_X2 _09429_ ( .A1(_02190_ ), .A2(_01805_ ), .A3(_02207_ ), .ZN(_02208_ ) );
NOR2_X1 _09430_ ( .A1(_02208_ ), .A2(_01833_ ), .ZN(_02209_ ) );
OR2_X1 _09431_ ( .A1(\ea_addr [11] ), .A2(ea_err ), .ZN(_02210_ ) );
OAI211_X1 _09432_ ( .A(_02129_ ), .B(_02210_ ), .C1(_00789_ ), .C2(\ea_pc [11] ), .ZN(_02211_ ) );
AND3_X1 _09433_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][11] ), .A3(_01579_ ), .ZN(_02212_ ) );
AND3_X1 _09434_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][11] ), .A3(_01462_ ), .ZN(_02213_ ) );
AOI21_X1 _09435_ ( .A(_02213_ ), .B1(_01584_ ), .B2(_01588_ ), .ZN(_02214_ ) );
NAND4_X1 _09436_ ( .A1(_01584_ ), .A2(\u_csr.csr[2][11] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_02215_ ) );
NAND2_X1 _09437_ ( .A1(_02214_ ), .A2(_02215_ ), .ZN(_02216_ ) );
OAI21_X1 _09438_ ( .A(_01576_ ), .B1(_02212_ ), .B2(_02216_ ), .ZN(_02217_ ) );
AND2_X1 _09439_ ( .A1(_02211_ ), .A2(_02217_ ), .ZN(_02218_ ) );
INV_X1 _09440_ ( .A(\de_pc [11] ), .ZN(_02219_ ) );
OAI22_X1 _09441_ ( .A1(_02218_ ), .A2(_01843_ ), .B1(_02219_ ), .B2(_01845_ ), .ZN(_02220_ ) );
OAI21_X1 _09442_ ( .A(_01855_ ), .B1(_02209_ ), .B2(_02220_ ), .ZN(_02221_ ) );
OAI22_X1 _09443_ ( .A1(_02208_ ), .A2(_01848_ ), .B1(_02219_ ), .B2(_01849_ ), .ZN(_02222_ ) );
AND3_X1 _09444_ ( .A1(_00672_ ), .A2(\u_idu.imm_branch [11] ), .A3(_00683_ ), .ZN(_02223_ ) );
AOI21_X1 _09445_ ( .A(_02223_ ), .B1(\u_idu.imm_auipc_lui [20] ), .B2(_00721_ ), .ZN(_02224_ ) );
OAI21_X1 _09446_ ( .A(_02224_ ), .B1(_00860_ ), .B2(_01091_ ), .ZN(_02225_ ) );
NOR2_X1 _09447_ ( .A1(_01780_ ), .A2(_02225_ ), .ZN(_02226_ ) );
INV_X1 _09448_ ( .A(_02226_ ), .ZN(_02227_ ) );
AOI21_X1 _09449_ ( .A(_02222_ ), .B1(_01495_ ), .B2(_02227_ ), .ZN(_02228_ ) );
OAI21_X1 _09450_ ( .A(_02221_ ), .B1(_02228_ ), .B2(_01854_ ), .ZN(_00142_ ) );
AND3_X1 _09451_ ( .A1(_01798_ ), .A2(_01143_ ), .A3(_01800_ ), .ZN(_02229_ ) );
AOI21_X1 _09452_ ( .A(_02229_ ), .B1(_02004_ ), .B2(_01796_ ), .ZN(_02230_ ) );
MUX2_X1 _09453_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ), .B(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ), .S(_01242_ ), .Z(_02231_ ) );
OAI21_X1 _09454_ ( .A(_01526_ ), .B1(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .B2(_02231_ ), .ZN(_02232_ ) );
OAI21_X1 _09455_ ( .A(_02232_ ), .B1(\io_master_rdata [10] ), .B2(_01526_ ), .ZN(_02233_ ) );
OAI21_X1 _09456_ ( .A(_02230_ ), .B1(_01277_ ), .B2(_02233_ ), .ZN(_02234_ ) );
AOI21_X2 _09457_ ( .A(_01604_ ), .B1(_01958_ ), .B2(_02234_ ), .ZN(_02235_ ) );
NAND2_X1 _09458_ ( .A1(_02235_ ), .A2(fanout_net_10 ), .ZN(_02236_ ) );
MUX2_X1 _09459_ ( .A(\u_exu.ecsr [10] ), .B(\ea_addr [10] ), .S(_01135_ ), .Z(_02237_ ) );
OR2_X1 _09460_ ( .A1(_02237_ ), .A2(fanout_net_10 ), .ZN(_02238_ ) );
AOI21_X1 _09461_ ( .A(_01686_ ), .B1(_02236_ ), .B2(_02238_ ), .ZN(_02239_ ) );
AOI22_X1 _09462_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02240_ ) );
AOI22_X1 _09463_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02241_ ) );
NAND3_X1 _09464_ ( .A1(_02240_ ), .A2(_01361_ ), .A3(_02241_ ), .ZN(_02242_ ) );
BUF_X4 _09465_ ( .A(_01336_ ), .Z(_02243_ ) );
OAI211_X1 _09466_ ( .A(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_02243_ ), .C1(_01871_ ), .C2(_01872_ ), .ZN(_02244_ ) );
INV_X1 _09467_ ( .A(\u_reg.rf[1][10] ), .ZN(_02245_ ) );
AOI21_X1 _09468_ ( .A(_01343_ ), .B1(_01345_ ), .B2(_02245_ ), .ZN(_02246_ ) );
NOR2_X1 _09469_ ( .A1(_01345_ ), .A2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02247_ ) );
OAI211_X1 _09470_ ( .A(_01335_ ), .B(_02244_ ), .C1(_02246_ ), .C2(_02247_ ), .ZN(_02248_ ) );
NAND3_X1 _09471_ ( .A1(_02242_ ), .A2(_01813_ ), .A3(_02248_ ), .ZN(_02249_ ) );
AOI22_X1 _09472_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02250_ ) );
AOI22_X1 _09473_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02251_ ) );
NAND3_X1 _09474_ ( .A1(_02250_ ), .A2(_01354_ ), .A3(_02251_ ), .ZN(_02252_ ) );
AOI22_X1 _09475_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02253_ ) );
AOI22_X1 _09476_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02254_ ) );
NAND3_X1 _09477_ ( .A1(_02253_ ), .A2(_01633_ ), .A3(_02254_ ), .ZN(_02255_ ) );
NAND3_X1 _09478_ ( .A1(_02252_ ), .A2(_02255_ ), .A3(_01705_ ), .ZN(_02256_ ) );
AOI21_X1 _09479_ ( .A(_01688_ ), .B1(_02249_ ), .B2(_02256_ ), .ZN(_02257_ ) );
NOR3_X2 _09480_ ( .A1(_02239_ ), .A2(_01317_ ), .A3(_02257_ ), .ZN(_02258_ ) );
NAND2_X1 _09481_ ( .A1(_02258_ ), .A2(_01370_ ), .ZN(_02259_ ) );
AND3_X1 _09482_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][10] ), .A3(_01461_ ), .ZN(_02260_ ) );
AOI21_X1 _09483_ ( .A(_02260_ ), .B1(_01588_ ), .B2(_01644_ ), .ZN(_02261_ ) );
NAND3_X1 _09484_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][10] ), .A3(_01647_ ), .ZN(_02262_ ) );
NAND4_X1 _09485_ ( .A1(_01651_ ), .A2(\u_csr.csr[2][10] ), .A3(_01648_ ), .A4(_01467_ ), .ZN(_02263_ ) );
NAND3_X1 _09486_ ( .A1(_02261_ ), .A2(_02262_ ), .A3(_02263_ ), .ZN(_02264_ ) );
NAND3_X1 _09487_ ( .A1(_01439_ ), .A2(_01444_ ), .A3(_02264_ ), .ZN(_02265_ ) );
NAND4_X1 _09488_ ( .A1(_01774_ ), .A2(_00813_ ), .A3(_00812_ ), .A4(_01715_ ), .ZN(_02266_ ) );
AOI21_X1 _09489_ ( .A(_01767_ ), .B1(_02265_ ), .B2(_02266_ ), .ZN(_02267_ ) );
AOI221_X4 _09490_ ( .A(_02267_ ), .B1(\de_pc [10] ), .B2(_01480_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_02268_ ) );
NAND2_X1 _09491_ ( .A1(_02258_ ), .A2(_01484_ ), .ZN(_02269_ ) );
AOI21_X1 _09492_ ( .A(_00861_ ), .B1(_01497_ ), .B2(_01832_ ), .ZN(_02270_ ) );
NOR3_X1 _09493_ ( .A1(_01779_ ), .A2(_00898_ ), .A3(\u_exu.opt_$_NOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B ), .ZN(_02271_ ) );
NOR2_X1 _09494_ ( .A1(_02270_ ), .A2(_02271_ ), .ZN(_02272_ ) );
INV_X1 _09495_ ( .A(_02272_ ), .ZN(_02273_ ) );
AOI221_X1 _09496_ ( .A(_01487_ ), .B1(\de_pc [10] ), .B2(_01491_ ), .C1(_01720_ ), .C2(_02273_ ), .ZN(_02274_ ) );
AOI221_X1 _09497_ ( .A(_00893_ ), .B1(_02259_ ), .B2(_02268_ ), .C1(_02269_ ), .C2(_02274_ ), .ZN(_00143_ ) );
BUF_X4 _09498_ ( .A(_00892_ ), .Z(_02275_ ) );
AND2_X1 _09499_ ( .A1(io_master_rready ), .A2(\io_master_rdata [9] ), .ZN(_02276_ ) );
MUX2_X1 _09500_ ( .A(\u_lsu.u_clint.mtime [41] ), .B(\u_lsu.u_clint.mtime [9] ), .S(_01529_ ), .Z(_02277_ ) );
AND3_X1 _09501_ ( .A1(_01527_ ), .A2(\u_lsu.rvalid_clint ), .A3(_02277_ ), .ZN(_02278_ ) );
NOR3_X1 _09502_ ( .A1(_02276_ ), .A2(_01276_ ), .A3(_02278_ ), .ZN(_02279_ ) );
AOI21_X1 _09503_ ( .A(_01144_ ), .B1(_01881_ ), .B2(_01882_ ), .ZN(_02280_ ) );
INV_X1 _09504_ ( .A(_01887_ ), .ZN(_02281_ ) );
AOI21_X1 _09505_ ( .A(_02280_ ), .B1(_02281_ ), .B2(_02004_ ), .ZN(_02282_ ) );
AOI211_X1 _09506_ ( .A(_01274_ ), .B(_02279_ ), .C1(_02282_ ), .C2(_01276_ ), .ZN(_02283_ ) );
OR3_X1 _09507_ ( .A1(_01604_ ), .A2(_01281_ ), .A3(_02283_ ), .ZN(_02284_ ) );
MUX2_X1 _09508_ ( .A(\u_exu.ecsr [9] ), .B(\ea_addr [9] ), .S(_01135_ ), .Z(_02285_ ) );
OR2_X1 _09509_ ( .A1(_02285_ ), .A2(fanout_net_10 ), .ZN(_02286_ ) );
AOI21_X1 _09510_ ( .A(_01312_ ), .B1(_02284_ ), .B2(_02286_ ), .ZN(_02287_ ) );
AOI22_X1 _09511_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02288_ ) );
AOI22_X1 _09512_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02289_ ) );
NAND3_X1 _09513_ ( .A1(_02288_ ), .A2(_01361_ ), .A3(_02289_ ), .ZN(_02290_ ) );
NAND3_X1 _09514_ ( .A1(_01546_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01338_ ), .ZN(_02291_ ) );
NOR2_X1 _09515_ ( .A1(_01551_ ), .A2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02292_ ) );
INV_X1 _09516_ ( .A(\u_reg.rf[1][9] ), .ZN(_02293_ ) );
AOI21_X1 _09517_ ( .A(_01694_ ), .B1(_01928_ ), .B2(_02293_ ), .ZN(_02294_ ) );
OAI211_X1 _09518_ ( .A(_02291_ ), .B(_01557_ ), .C1(_02292_ ), .C2(_02294_ ), .ZN(_02295_ ) );
NAND3_X1 _09519_ ( .A1(_02290_ ), .A2(_01813_ ), .A3(_02295_ ), .ZN(_02296_ ) );
AOI22_X1 _09520_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02297_ ) );
AOI22_X1 _09521_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02298_ ) );
NAND3_X1 _09522_ ( .A1(_02297_ ), .A2(_01335_ ), .A3(_02298_ ), .ZN(_02299_ ) );
AOI22_X1 _09523_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02300_ ) );
AOI22_X1 _09524_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02301_ ) );
NAND3_X1 _09525_ ( .A1(_02300_ ), .A2(_01633_ ), .A3(_02301_ ), .ZN(_02302_ ) );
NAND3_X1 _09526_ ( .A1(_02299_ ), .A2(_02302_ ), .A3(_01705_ ), .ZN(_02303_ ) );
AOI21_X1 _09527_ ( .A(_01688_ ), .B1(_02296_ ), .B2(_02303_ ), .ZN(_02304_ ) );
NOR3_X2 _09528_ ( .A1(_02287_ ), .A2(_01316_ ), .A3(_02304_ ), .ZN(_02305_ ) );
NAND2_X1 _09529_ ( .A1(_02305_ ), .A2(_01370_ ), .ZN(_02306_ ) );
AND3_X1 _09530_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][9] ), .A3(_01647_ ), .ZN(_02307_ ) );
NAND4_X1 _09531_ ( .A1(_01582_ ), .A2(\u_csr.csr[2][9] ), .A3(_00754_ ), .A4(_01591_ ), .ZN(_02308_ ) );
NAND3_X1 _09532_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][9] ), .A3(_01461_ ), .ZN(_02309_ ) );
NAND2_X1 _09533_ ( .A1(_02308_ ), .A2(_02309_ ), .ZN(_02310_ ) );
OAI21_X1 _09534_ ( .A(_01575_ ), .B1(_02307_ ), .B2(_02310_ ), .ZN(_02311_ ) );
NAND4_X1 _09535_ ( .A1(_01774_ ), .A2(_00817_ ), .A3(_00816_ ), .A4(_01715_ ), .ZN(_02312_ ) );
AOI21_X1 _09536_ ( .A(_01767_ ), .B1(_02311_ ), .B2(_02312_ ), .ZN(_02313_ ) );
AOI221_X4 _09537_ ( .A(_02313_ ), .B1(\de_pc [9] ), .B2(_01480_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_02314_ ) );
NAND2_X1 _09538_ ( .A1(_02305_ ), .A2(_01484_ ), .ZN(_02315_ ) );
AOI21_X1 _09539_ ( .A(_00881_ ), .B1(_01497_ ), .B2(_01514_ ), .ZN(_02316_ ) );
AOI221_X1 _09540_ ( .A(_01487_ ), .B1(\de_pc [9] ), .B2(_01491_ ), .C1(_01720_ ), .C2(_02316_ ), .ZN(_02317_ ) );
AOI221_X1 _09541_ ( .A(_02275_ ), .B1(_02306_ ), .B2(_02314_ ), .C1(_02315_ ), .C2(_02317_ ), .ZN(_00144_ ) );
AND3_X1 _09542_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [8] ), .ZN(_02318_ ) );
AOI211_X1 _09543_ ( .A(fanout_net_10 ), .B(_02318_ ), .C1(\ea_addr [8] ), .C2(_01521_ ), .ZN(_02319_ ) );
AND3_X1 _09544_ ( .A1(_01914_ ), .A2(_01143_ ), .A3(_01918_ ), .ZN(_02320_ ) );
AOI21_X1 _09545_ ( .A(_02320_ ), .B1(_02004_ ), .B2(_01912_ ), .ZN(_02321_ ) );
MUX2_X1 _09546_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ), .B(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ), .S(_01529_ ), .Z(_02322_ ) );
OAI21_X1 _09547_ ( .A(_01527_ ), .B1(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .B2(_02322_ ), .ZN(_02323_ ) );
OAI21_X1 _09548_ ( .A(_02323_ ), .B1(\io_master_rdata [8] ), .B2(_01909_ ), .ZN(_02324_ ) );
OAI21_X1 _09549_ ( .A(_02321_ ), .B1(_01277_ ), .B2(_02324_ ), .ZN(_02325_ ) );
AOI21_X2 _09550_ ( .A(_01604_ ), .B1(_01958_ ), .B2(_02325_ ), .ZN(_02326_ ) );
AOI21_X2 _09551_ ( .A(_02319_ ), .B1(_02326_ ), .B2(fanout_net_10 ), .ZN(\ar_data [8] ) );
NOR2_X1 _09552_ ( .A1(\ar_data [8] ), .A2(_01313_ ), .ZN(_02327_ ) );
AOI22_X1 _09553_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02328_ ) );
AOI22_X1 _09554_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02329_ ) );
NAND3_X1 _09555_ ( .A1(_02328_ ), .A2(_01809_ ), .A3(_02329_ ), .ZN(_02330_ ) );
NAND3_X1 _09556_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01547_ ), .ZN(_02331_ ) );
NOR2_X1 _09557_ ( .A1(_01549_ ), .A2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02332_ ) );
INV_X1 _09558_ ( .A(\u_reg.rf[1][8] ), .ZN(_02333_ ) );
AOI21_X1 _09559_ ( .A(_01343_ ), .B1(_01551_ ), .B2(_02333_ ), .ZN(_02334_ ) );
OAI211_X1 _09560_ ( .A(_02331_ ), .B(_01558_ ), .C1(_02332_ ), .C2(_02334_ ), .ZN(_02335_ ) );
NAND3_X1 _09561_ ( .A1(_02330_ ), .A2(_01814_ ), .A3(_02335_ ), .ZN(_02336_ ) );
AOI22_X1 _09562_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02337_ ) );
AOI22_X1 _09563_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02338_ ) );
AOI21_X1 _09564_ ( .A(_01354_ ), .B1(_02337_ ), .B2(_02338_ ), .ZN(_02339_ ) );
AOI22_X1 _09565_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01322_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02340_ ) );
AOI22_X1 _09566_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02341_ ) );
AOI21_X1 _09567_ ( .A(_01361_ ), .B1(_02340_ ), .B2(_02341_ ), .ZN(_02342_ ) );
OAI21_X1 _09568_ ( .A(_01822_ ), .B1(_02339_ ), .B2(_02342_ ), .ZN(_02343_ ) );
AOI21_X1 _09569_ ( .A(_01318_ ), .B1(_02336_ ), .B2(_02343_ ), .ZN(_02344_ ) );
OR3_X2 _09570_ ( .A1(_02327_ ), .A2(_01317_ ), .A3(_02344_ ), .ZN(_02345_ ) );
NOR2_X1 _09571_ ( .A1(_02345_ ), .A2(_01833_ ), .ZN(_02346_ ) );
AND3_X1 _09572_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][8] ), .A3(_01579_ ), .ZN(_02347_ ) );
AND3_X1 _09573_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][8] ), .A3(_01462_ ), .ZN(_02348_ ) );
AOI21_X1 _09574_ ( .A(_02348_ ), .B1(_01583_ ), .B2(_01588_ ), .ZN(_02349_ ) );
NAND4_X1 _09575_ ( .A1(_01583_ ), .A2(\u_csr.csr[2][8] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_02350_ ) );
NAND2_X1 _09576_ ( .A1(_02349_ ), .A2(_02350_ ), .ZN(_02351_ ) );
OAI21_X1 _09577_ ( .A(_01576_ ), .B1(_02347_ ), .B2(_02351_ ), .ZN(_02352_ ) );
NAND4_X1 _09578_ ( .A1(_01596_ ), .A2(_00819_ ), .A3(_00818_ ), .A4(_01444_ ), .ZN(_02353_ ) );
AND2_X1 _09579_ ( .A1(_02352_ ), .A2(_02353_ ), .ZN(_02354_ ) );
INV_X1 _09580_ ( .A(\de_pc [8] ), .ZN(_02355_ ) );
OAI22_X1 _09581_ ( .A1(_02354_ ), .A2(_01843_ ), .B1(_02355_ ), .B2(_01845_ ), .ZN(_02356_ ) );
OAI21_X1 _09582_ ( .A(_01855_ ), .B1(_02346_ ), .B2(_02356_ ), .ZN(_02357_ ) );
OAI22_X1 _09583_ ( .A1(_02345_ ), .A2(_01483_ ), .B1(_02355_ ), .B2(_01849_ ), .ZN(_02358_ ) );
AND2_X2 _09584_ ( .A1(_01497_ ), .A2(_01514_ ), .ZN(_02359_ ) );
NOR2_X1 _09585_ ( .A1(_02359_ ), .A2(_00884_ ), .ZN(_02360_ ) );
AOI21_X1 _09586_ ( .A(_02358_ ), .B1(_01495_ ), .B2(_02360_ ), .ZN(_02361_ ) );
OAI21_X1 _09587_ ( .A(_02357_ ), .B1(_02361_ ), .B2(_01570_ ), .ZN(_00145_ ) );
BUF_X4 _09588_ ( .A(_01490_ ), .Z(_02362_ ) );
NAND3_X1 _09589_ ( .A1(_01483_ ), .A2(\de_pc [7] ), .A3(_02362_ ), .ZN(_02363_ ) );
MUX2_X1 _09590_ ( .A(\u_exu.ecsr [7] ), .B(\ea_addr [7] ), .S(_01135_ ), .Z(_02364_ ) );
AND2_X1 _09591_ ( .A1(_01260_ ), .A2(_01270_ ), .ZN(_02365_ ) );
NOR2_X1 _09592_ ( .A1(_01259_ ), .A2(_02365_ ), .ZN(_02366_ ) );
MUX2_X1 _09593_ ( .A(_02364_ ), .B(_02366_ ), .S(fanout_net_10 ), .Z(\ar_data [7] ) );
NOR2_X1 _09594_ ( .A1(\ar_data [7] ), .A2(_01686_ ), .ZN(_02367_ ) );
AOI22_X1 _09595_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02368_ ) );
AOI22_X1 _09596_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02369_ ) );
NAND3_X1 _09597_ ( .A1(_02368_ ), .A2(_01633_ ), .A3(_02369_ ), .ZN(_02370_ ) );
OAI211_X1 _09598_ ( .A(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_02243_ ), .C1(_01871_ ), .C2(_01872_ ), .ZN(_02371_ ) );
INV_X1 _09599_ ( .A(\u_reg.rf[1][7] ), .ZN(_02372_ ) );
AOI21_X1 _09600_ ( .A(_01694_ ), .B1(_01928_ ), .B2(_02372_ ), .ZN(_02373_ ) );
NOR2_X1 _09601_ ( .A1(_01928_ ), .A2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02374_ ) );
OAI211_X1 _09602_ ( .A(_01557_ ), .B(_02371_ ), .C1(_02373_ ), .C2(_02374_ ), .ZN(_02375_ ) );
NAND3_X1 _09603_ ( .A1(_02370_ ), .A2(_01813_ ), .A3(_02375_ ), .ZN(_02376_ ) );
AOI22_X1 _09604_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02377_ ) );
AOI22_X1 _09605_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01752_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02378_ ) );
NAND3_X1 _09606_ ( .A1(_02377_ ), .A2(_01335_ ), .A3(_02378_ ), .ZN(_02379_ ) );
AOI22_X1 _09607_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02380_ ) );
AOI22_X1 _09608_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01752_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02381_ ) );
NAND3_X1 _09609_ ( .A1(_02380_ ), .A2(_01756_ ), .A3(_02381_ ), .ZN(_02382_ ) );
NAND3_X1 _09610_ ( .A1(_02379_ ), .A2(_02382_ ), .A3(_01705_ ), .ZN(_02383_ ) );
AOI21_X2 _09611_ ( .A(_01688_ ), .B1(_02376_ ), .B2(_02383_ ), .ZN(_02384_ ) );
OR3_X2 _09612_ ( .A1(_02367_ ), .A2(_01316_ ), .A3(_02384_ ), .ZN(_02385_ ) );
OAI21_X1 _09613_ ( .A(_02363_ ), .B1(_02385_ ), .B2(_01848_ ), .ZN(_02386_ ) );
NOR2_X1 _09614_ ( .A1(_02359_ ), .A2(_00886_ ), .ZN(_02387_ ) );
AND3_X1 _09615_ ( .A1(_00709_ ), .A2(_01493_ ), .A3(_02387_ ), .ZN(_02388_ ) );
OAI21_X1 _09616_ ( .A(_01569_ ), .B1(_02386_ ), .B2(_02388_ ), .ZN(_02389_ ) );
OR2_X2 _09617_ ( .A1(_02385_ ), .A2(_01832_ ), .ZN(_02390_ ) );
AND3_X1 _09618_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][7] ), .A3(_01579_ ), .ZN(_02391_ ) );
NAND4_X1 _09619_ ( .A1(_01583_ ), .A2(\u_csr.csr[2][7] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_02392_ ) );
AND3_X1 _09620_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][7] ), .A3(_01462_ ), .ZN(_02393_ ) );
AOI21_X1 _09621_ ( .A(_02393_ ), .B1(_01588_ ), .B2(_01644_ ), .ZN(_02394_ ) );
NAND2_X1 _09622_ ( .A1(_02392_ ), .A2(_02394_ ), .ZN(_02395_ ) );
OAI21_X1 _09623_ ( .A(_01576_ ), .B1(_02391_ ), .B2(_02395_ ), .ZN(_02396_ ) );
NAND4_X1 _09624_ ( .A1(_01596_ ), .A2(_00821_ ), .A3(_00820_ ), .A4(_01597_ ), .ZN(_02397_ ) );
AND2_X1 _09625_ ( .A1(_02396_ ), .A2(_02397_ ), .ZN(_02398_ ) );
OR2_X1 _09626_ ( .A1(_02398_ ), .A2(_01375_ ), .ZN(_02399_ ) );
OAI21_X1 _09627_ ( .A(\de_pc [7] ), .B1(_01476_ ), .B2(_01477_ ), .ZN(_02400_ ) );
AND3_X2 _09628_ ( .A1(_02390_ ), .A2(_02399_ ), .A3(_02400_ ), .ZN(_02401_ ) );
OAI21_X1 _09629_ ( .A(_02389_ ), .B1(_02401_ ), .B2(_01572_ ), .ZN(_00146_ ) );
INV_X1 _09630_ ( .A(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02402_ ) );
INV_X1 _09631_ ( .A(_01017_ ), .ZN(_02403_ ) );
INV_X1 _09632_ ( .A(_01321_ ), .ZN(_02404_ ) );
INV_X1 _09633_ ( .A(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02405_ ) );
OAI22_X1 _09634_ ( .A1(_02402_ ), .A2(_02403_ ), .B1(_02404_ ), .B2(_02405_ ), .ZN(_02406_ ) );
OAI211_X1 _09635_ ( .A(_01342_ ), .B(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C1(_00933_ ), .C2(_00934_ ), .ZN(_02407_ ) );
INV_X1 _09636_ ( .A(_01329_ ), .ZN(_02408_ ) );
INV_X1 _09637_ ( .A(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02409_ ) );
OAI21_X1 _09638_ ( .A(_02407_ ), .B1(_02408_ ), .B2(_02409_ ), .ZN(_02410_ ) );
OAI21_X1 _09639_ ( .A(_01756_ ), .B1(_02406_ ), .B2(_02410_ ), .ZN(_02411_ ) );
AOI22_X1 _09640_ ( .A1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01327_ ), .B1(_01330_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02412_ ) );
NAND3_X1 _09641_ ( .A1(_01344_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01342_ ), .ZN(_02413_ ) );
NAND3_X1 _09642_ ( .A1(_01344_ ), .A2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01337_ ), .ZN(_02414_ ) );
AND3_X1 _09643_ ( .A1(_02412_ ), .A2(_02413_ ), .A3(_02414_ ), .ZN(_02415_ ) );
OAI211_X1 _09644_ ( .A(_02411_ ), .B(_01705_ ), .C1(_01326_ ), .C2(_02415_ ), .ZN(_02416_ ) );
MUX2_X1 _09645_ ( .A(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_01336_ ), .Z(_02417_ ) );
AND2_X1 _09646_ ( .A1(_02417_ ), .A2(_01344_ ), .ZN(_02418_ ) );
OAI211_X1 _09647_ ( .A(_01342_ ), .B(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C1(_00933_ ), .C2(_00934_ ), .ZN(_02419_ ) );
OAI211_X1 _09648_ ( .A(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(_01337_ ), .C1(_00933_ ), .C2(_00934_ ), .ZN(_02420_ ) );
NAND2_X1 _09649_ ( .A1(_02419_ ), .A2(_02420_ ), .ZN(_02421_ ) );
OAI21_X1 _09650_ ( .A(_01756_ ), .B1(_02418_ ), .B2(_02421_ ), .ZN(_02422_ ) );
OAI21_X1 _09651_ ( .A(_01342_ ), .B1(_01344_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02423_ ) );
OAI21_X1 _09652_ ( .A(_02423_ ), .B1(\u_reg.rf[1][6] ), .B2(_01545_ ), .ZN(_02424_ ) );
AOI21_X1 _09653_ ( .A(_02424_ ), .B1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_01810_ ), .ZN(_02425_ ) );
OAI211_X1 _09654_ ( .A(_02422_ ), .B(_01813_ ), .C1(_02425_ ), .C2(_01326_ ), .ZN(_02426_ ) );
AND3_X1 _09655_ ( .A1(_01312_ ), .A2(_02416_ ), .A3(_02426_ ), .ZN(_02427_ ) );
MUX2_X1 _09656_ ( .A(\u_exu.ecsr [6] ), .B(\ea_addr [6] ), .S(_01135_ ), .Z(_02428_ ) );
NOR2_X1 _09657_ ( .A1(_02428_ ), .A2(fanout_net_10 ), .ZN(_02429_ ) );
INV_X1 _09658_ ( .A(_02365_ ), .ZN(_02430_ ) );
BUF_X2 _09659_ ( .A(_02430_ ), .Z(_02431_ ) );
AND3_X1 _09660_ ( .A1(_01998_ ), .A2(_02004_ ), .A3(_02002_ ), .ZN(_02432_ ) );
AOI21_X1 _09661_ ( .A(_02432_ ), .B1(_01236_ ), .B2(_01532_ ), .ZN(_02433_ ) );
OAI21_X1 _09662_ ( .A(_02433_ ), .B1(_01144_ ), .B2(_02008_ ), .ZN(_02434_ ) );
MUX2_X1 _09663_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ), .B(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ), .S(_01733_ ), .Z(_02435_ ) );
OR4_X1 _09664_ ( .A1(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .A2(_01607_ ), .A3(_01608_ ), .A4(_02435_ ), .ZN(_02436_ ) );
OAI21_X1 _09665_ ( .A(\io_master_rdata [6] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_02437_ ) );
AOI21_X1 _09666_ ( .A(_01277_ ), .B1(_02436_ ), .B2(_02437_ ), .ZN(_02438_ ) );
OAI21_X1 _09667_ ( .A(_02431_ ), .B1(_02434_ ), .B2(_02438_ ), .ZN(_02439_ ) );
AOI21_X2 _09668_ ( .A(_02429_ ), .B1(_02439_ ), .B2(fanout_net_10 ), .ZN(\ar_data [6] ) );
NOR2_X1 _09669_ ( .A1(\ar_data [6] ), .A2(_01686_ ), .ZN(_02440_ ) );
NOR3_X2 _09670_ ( .A1(_02427_ ), .A2(_02440_ ), .A3(_01316_ ), .ZN(_02441_ ) );
NAND2_X1 _09671_ ( .A1(_02441_ ), .A2(_01370_ ), .ZN(_02442_ ) );
NAND4_X1 _09672_ ( .A1(_01455_ ), .A2(\u_csr.csr[2][6] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_02443_ ) );
NAND3_X1 _09673_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][6] ), .A3(_01647_ ), .ZN(_02444_ ) );
NAND4_X1 _09674_ ( .A1(_01653_ ), .A2(\u_csr.csr[0][6] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_02445_ ) );
NAND4_X1 _09675_ ( .A1(_01646_ ), .A2(_02443_ ), .A3(_02444_ ), .A4(_02445_ ), .ZN(_02446_ ) );
NAND2_X1 _09676_ ( .A1(_01576_ ), .A2(_02446_ ), .ZN(_02447_ ) );
NAND4_X1 _09677_ ( .A1(_01774_ ), .A2(_00823_ ), .A3(_00822_ ), .A4(_01715_ ), .ZN(_02448_ ) );
AOI21_X1 _09678_ ( .A(_01767_ ), .B1(_02447_ ), .B2(_02448_ ), .ZN(_02449_ ) );
AOI221_X4 _09679_ ( .A(_02449_ ), .B1(\de_pc [6] ), .B2(_01479_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_02450_ ) );
NAND2_X1 _09680_ ( .A1(_02441_ ), .A2(_01484_ ), .ZN(_02451_ ) );
NOR2_X1 _09681_ ( .A1(_02359_ ), .A2(_00732_ ), .ZN(_02452_ ) );
AOI221_X1 _09682_ ( .A(_01487_ ), .B1(\de_pc [6] ), .B2(_01491_ ), .C1(_01720_ ), .C2(_02452_ ), .ZN(_02453_ ) );
AOI221_X1 _09683_ ( .A(_02275_ ), .B1(_02442_ ), .B2(_02450_ ), .C1(_02451_ ), .C2(_02453_ ), .ZN(_00147_ ) );
BUF_X4 _09684_ ( .A(_00892_ ), .Z(_02454_ ) );
BUF_X4 _09685_ ( .A(_02454_ ), .Z(_02455_ ) );
BUF_X4 _09686_ ( .A(_02455_ ), .Z(_02456_ ) );
AOI21_X1 _09687_ ( .A(_00656_ ), .B1(_01497_ ), .B2(_01514_ ), .ZN(_02457_ ) );
NAND3_X1 _09688_ ( .A1(_00709_ ), .A2(_01493_ ), .A3(_02457_ ), .ZN(_02458_ ) );
INV_X1 _09689_ ( .A(\de_pc [5] ), .ZN(_02459_ ) );
MUX2_X1 _09690_ ( .A(\u_exu.ecsr [5] ), .B(\ea_addr [5] ), .S(_01136_ ), .Z(_02460_ ) );
OAI21_X1 _09691_ ( .A(_01143_ ), .B1(_02057_ ), .B2(_02058_ ), .ZN(_02461_ ) );
OAI21_X1 _09692_ ( .A(_02461_ ), .B1(_01610_ ), .B2(_01247_ ), .ZN(_02462_ ) );
AOI21_X1 _09693_ ( .A(_01237_ ), .B1(_01612_ ), .B2(_01613_ ), .ZN(_02463_ ) );
OR3_X2 _09694_ ( .A1(_02462_ ), .A2(_01524_ ), .A3(_02463_ ), .ZN(_02464_ ) );
AOI21_X1 _09695_ ( .A(_01276_ ), .B1(io_master_rready ), .B2(\io_master_rdata [5] ), .ZN(_02465_ ) );
AND3_X1 _09696_ ( .A1(_01669_ ), .A2(\u_lsu.u_clint.mtime [5] ), .A3(_01524_ ), .ZN(_02466_ ) );
AOI21_X1 _09697_ ( .A(_02466_ ), .B1(_01249_ ), .B2(\u_lsu.u_clint.mtime [37] ), .ZN(_02467_ ) );
OAI21_X1 _09698_ ( .A(_02465_ ), .B1(_01229_ ), .B2(_02467_ ), .ZN(_02468_ ) );
AND3_X2 _09699_ ( .A1(_02464_ ), .A2(_02431_ ), .A3(_02468_ ), .ZN(_02469_ ) );
MUX2_X2 _09700_ ( .A(_02460_ ), .B(_02469_ ), .S(fanout_net_10 ), .Z(\ar_data [5] ) );
AND2_X2 _09701_ ( .A1(\ar_data [5] ), .A2(_01318_ ), .ZN(_02470_ ) );
AOI22_X1 _09702_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_02012_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02471_ ) );
AOI22_X1 _09703_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02472_ ) );
NAND3_X1 _09704_ ( .A1(_02471_ ), .A2(_02015_ ), .A3(_02472_ ), .ZN(_02473_ ) );
NAND3_X1 _09705_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01965_ ), .ZN(_02474_ ) );
NOR2_X1 _09706_ ( .A1(_02021_ ), .A2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02475_ ) );
INV_X1 _09707_ ( .A(\u_reg.rf[1][5] ), .ZN(_02476_ ) );
AOI21_X1 _09708_ ( .A(_01816_ ), .B1(_02021_ ), .B2(_02476_ ), .ZN(_02477_ ) );
OAI211_X1 _09709_ ( .A(_02474_ ), .B(_01858_ ), .C1(_02475_ ), .C2(_02477_ ), .ZN(_02478_ ) );
NAND3_X1 _09710_ ( .A1(_02473_ ), .A2(_01814_ ), .A3(_02478_ ), .ZN(_02479_ ) );
AOI22_X1 _09711_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_02012_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02480_ ) );
AOI22_X1 _09712_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02481_ ) );
AOI21_X1 _09713_ ( .A(_01858_ ), .B1(_02480_ ), .B2(_02481_ ), .ZN(_02482_ ) );
AOI22_X1 _09714_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02483_ ) );
AOI22_X1 _09715_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02484_ ) );
AOI21_X1 _09716_ ( .A(_01809_ ), .B1(_02483_ ), .B2(_02484_ ), .ZN(_02485_ ) );
OAI21_X1 _09717_ ( .A(_01822_ ), .B1(_02482_ ), .B2(_02485_ ), .ZN(_02486_ ) );
AND3_X1 _09718_ ( .A1(_01536_ ), .A2(_02479_ ), .A3(_02486_ ), .ZN(_02487_ ) );
OAI21_X1 _09719_ ( .A(_01535_ ), .B1(_02470_ ), .B2(_02487_ ), .ZN(_02488_ ) );
OAI221_X1 _09720_ ( .A(_02458_ ), .B1(_02459_ ), .B2(_01849_ ), .C1(_02488_ ), .C2(_01848_ ), .ZN(_02489_ ) );
NAND2_X1 _09721_ ( .A1(_02489_ ), .A2(_01090_ ), .ZN(_02490_ ) );
NOR2_X1 _09722_ ( .A1(_02488_ ), .A2(_01832_ ), .ZN(_02491_ ) );
INV_X4 _09723_ ( .A(_01574_ ), .ZN(_02492_ ) );
AND4_X1 _09724_ ( .A1(\u_csr.csr[0][5] ), .A2(_01653_ ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_02493_ ) );
AND2_X1 _09725_ ( .A1(_01450_ ), .A2(_01453_ ), .ZN(_02494_ ) );
AOI21_X1 _09726_ ( .A(_02493_ ), .B1(_02494_ ), .B2(\u_csr.csr[1][5] ), .ZN(_02495_ ) );
AND3_X1 _09727_ ( .A1(_01455_ ), .A2(_01590_ ), .A3(_01653_ ), .ZN(_02496_ ) );
AND3_X1 _09728_ ( .A1(_02496_ ), .A2(\u_csr.csr[2][5] ), .A3(_01592_ ), .ZN(_02497_ ) );
NOR3_X1 _09729_ ( .A1(_02497_ ), .A2(_01641_ ), .A3(_01645_ ), .ZN(_02498_ ) );
AOI21_X1 _09730_ ( .A(_02492_ ), .B1(_02495_ ), .B2(_02498_ ), .ZN(_02499_ ) );
NAND2_X1 _09731_ ( .A1(_00824_ ), .A2(_00825_ ), .ZN(_02500_ ) );
NAND4_X1 _09732_ ( .A1(_01398_ ), .A2(_01428_ ), .A3(_01379_ ), .A4(_01383_ ), .ZN(_02501_ ) );
NAND4_X1 _09733_ ( .A1(_01435_ ), .A2(_01386_ ), .A3(_01429_ ), .A4(_01436_ ), .ZN(_02502_ ) );
AND4_X1 _09734_ ( .A1(_01401_ ), .A2(_01400_ ), .A3(_01402_ ), .A4(_01415_ ), .ZN(_02503_ ) );
INV_X1 _09735_ ( .A(_01417_ ), .ZN(_02504_ ) );
INV_X1 _09736_ ( .A(_01416_ ), .ZN(_02505_ ) );
AND4_X1 _09737_ ( .A1(_02504_ ), .A2(_01412_ ), .A3(_02505_ ), .A4(_01408_ ), .ZN(_02506_ ) );
NAND2_X1 _09738_ ( .A1(_02503_ ), .A2(_02506_ ), .ZN(_02507_ ) );
NAND4_X1 _09739_ ( .A1(_01423_ ), .A2(_01432_ ), .A3(_01389_ ), .A4(_01421_ ), .ZN(_02508_ ) );
NOR4_X1 _09740_ ( .A1(_02501_ ), .A2(_02502_ ), .A3(_02507_ ), .A4(_02508_ ), .ZN(_02509_ ) );
AND4_X1 _09741_ ( .A1(_02500_ ), .A2(_02509_ ), .A3(_01597_ ), .A4(_01381_ ), .ZN(_02510_ ) );
OAI21_X1 _09742_ ( .A(_01373_ ), .B1(_02499_ ), .B2(_02510_ ), .ZN(_02511_ ) );
OAI21_X1 _09743_ ( .A(_02511_ ), .B1(_02459_ ), .B2(_01845_ ), .ZN(_02512_ ) );
OAI21_X1 _09744_ ( .A(_01057_ ), .B1(_02491_ ), .B2(_02512_ ), .ZN(_02513_ ) );
AOI21_X1 _09745_ ( .A(_02456_ ), .B1(_02490_ ), .B2(_02513_ ), .ZN(_00148_ ) );
MUX2_X1 _09746_ ( .A(\u_exu.ecsr [4] ), .B(\ea_addr [4] ), .S(_01136_ ), .Z(_02514_ ) );
AND3_X1 _09747_ ( .A1(_01678_ ), .A2(_02004_ ), .A3(_01682_ ), .ZN(_02515_ ) );
AOI21_X1 _09748_ ( .A(_02515_ ), .B1(_01236_ ), .B2(_01675_ ), .ZN(_02516_ ) );
NOR2_X1 _09749_ ( .A1(_02105_ ), .A2(_01144_ ), .ZN(_02517_ ) );
INV_X1 _09750_ ( .A(_02517_ ), .ZN(_02518_ ) );
AND3_X1 _09751_ ( .A1(_02516_ ), .A2(_01277_ ), .A3(_02518_ ), .ZN(_02519_ ) );
AND2_X1 _09752_ ( .A1(io_master_rready ), .A2(\io_master_rdata [4] ), .ZN(_02520_ ) );
AND3_X1 _09753_ ( .A1(_01669_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ), .A3(_01524_ ), .ZN(_02521_ ) );
INV_X1 _09754_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_26_A_$_ANDNOT__Y_B ), .ZN(_02522_ ) );
AOI21_X1 _09755_ ( .A(_02522_ ), .B1(_01669_ ), .B2(_01524_ ), .ZN(_02523_ ) );
NOR3_X1 _09756_ ( .A1(_02521_ ), .A2(_02523_ ), .A3(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .ZN(_02524_ ) );
AND2_X1 _09757_ ( .A1(_01909_ ), .A2(_02524_ ), .ZN(_02525_ ) );
NOR3_X1 _09758_ ( .A1(_02520_ ), .A2(_01277_ ), .A3(_02525_ ), .ZN(_02526_ ) );
NOR3_X1 _09759_ ( .A1(_02519_ ), .A2(_02365_ ), .A3(_02526_ ), .ZN(_02527_ ) );
MUX2_X2 _09760_ ( .A(_02514_ ), .B(_02527_ ), .S(fanout_net_10 ), .Z(\ar_data [4] ) );
NOR2_X1 _09761_ ( .A1(\ar_data [4] ), .A2(_01536_ ), .ZN(_02528_ ) );
AOI22_X1 _09762_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02529_ ) );
AOI22_X1 _09763_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02530_ ) );
AOI21_X1 _09764_ ( .A(_01325_ ), .B1(_02529_ ), .B2(_02530_ ), .ZN(_02531_ ) );
AOI22_X1 _09765_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01319_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02532_ ) );
AOI22_X1 _09766_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01330_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02533_ ) );
AOI21_X1 _09767_ ( .A(_01557_ ), .B1(_02532_ ), .B2(_02533_ ), .ZN(_02534_ ) );
OR3_X1 _09768_ ( .A1(_02531_ ), .A2(_02534_ ), .A3(_01813_ ), .ZN(_02535_ ) );
NAND3_X1 _09769_ ( .A1(_01928_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_02243_ ), .ZN(_02536_ ) );
INV_X1 _09770_ ( .A(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02537_ ) );
OAI21_X1 _09771_ ( .A(_02536_ ), .B1(_02403_ ), .B2(_02537_ ), .ZN(_02538_ ) );
OAI211_X1 _09772_ ( .A(_01694_ ), .B(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C1(_01871_ ), .C2(_01872_ ), .ZN(_02539_ ) );
OAI211_X1 _09773_ ( .A(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(_02243_ ), .C1(_01871_ ), .C2(_01872_ ), .ZN(_02540_ ) );
NAND2_X1 _09774_ ( .A1(_02539_ ), .A2(_02540_ ), .ZN(_02541_ ) );
OAI21_X1 _09775_ ( .A(_01326_ ), .B1(_02538_ ), .B2(_02541_ ), .ZN(_02542_ ) );
AND3_X1 _09776_ ( .A1(_01545_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_02243_ ), .ZN(_02543_ ) );
OR2_X1 _09777_ ( .A1(_01928_ ), .A2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02544_ ) );
OAI21_X1 _09778_ ( .A(_01547_ ), .B1(_01546_ ), .B2(\u_reg.rf[1][4] ), .ZN(_02545_ ) );
AOI21_X1 _09779_ ( .A(_02543_ ), .B1(_02544_ ), .B2(_02545_ ), .ZN(_02546_ ) );
OAI211_X1 _09780_ ( .A(_02542_ ), .B(_01334_ ), .C1(_02015_ ), .C2(_02546_ ), .ZN(_02547_ ) );
AND3_X2 _09781_ ( .A1(_01313_ ), .A2(_02535_ ), .A3(_02547_ ), .ZN(_02548_ ) );
NOR3_X1 _09782_ ( .A1(_02528_ ), .A2(_01805_ ), .A3(_02548_ ), .ZN(_02549_ ) );
AND2_X1 _09783_ ( .A1(_02549_ ), .A2(_01371_ ), .ZN(_02550_ ) );
AND3_X1 _09784_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][4] ), .A3(_01579_ ), .ZN(_02551_ ) );
AND3_X1 _09785_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][4] ), .A3(_01462_ ), .ZN(_02552_ ) );
AOI21_X1 _09786_ ( .A(_02552_ ), .B1(_01584_ ), .B2(_01588_ ), .ZN(_02553_ ) );
NAND4_X1 _09787_ ( .A1(_01584_ ), .A2(\u_csr.csr[2][4] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_02554_ ) );
NAND2_X1 _09788_ ( .A1(_02553_ ), .A2(_02554_ ), .ZN(_02555_ ) );
OAI21_X1 _09789_ ( .A(_01576_ ), .B1(_02551_ ), .B2(_02555_ ), .ZN(_02556_ ) );
NAND4_X1 _09790_ ( .A1(_01596_ ), .A2(_00827_ ), .A3(_00826_ ), .A4(_01597_ ), .ZN(_02557_ ) );
AND2_X1 _09791_ ( .A1(_02556_ ), .A2(_02557_ ), .ZN(_02558_ ) );
INV_X1 _09792_ ( .A(\de_pc [4] ), .ZN(_02559_ ) );
OAI22_X1 _09793_ ( .A1(_02558_ ), .A2(_01843_ ), .B1(_02559_ ), .B2(_01478_ ), .ZN(_02560_ ) );
OAI21_X1 _09794_ ( .A(_01855_ ), .B1(_02550_ ), .B2(_02560_ ), .ZN(_02561_ ) );
NAND2_X1 _09795_ ( .A1(_02549_ ), .A2(_01485_ ), .ZN(_02562_ ) );
INV_X1 _09796_ ( .A(_01496_ ), .ZN(_02563_ ) );
AND2_X1 _09797_ ( .A1(_02563_ ), .A2(\u_idu.imm_branch [4] ), .ZN(_02564_ ) );
AOI21_X1 _09798_ ( .A(_00887_ ), .B1(_00727_ ), .B2(_00895_ ), .ZN(_02565_ ) );
OR2_X1 _09799_ ( .A1(_02564_ ), .A2(_02565_ ), .ZN(_02566_ ) );
NAND3_X1 _09800_ ( .A1(_00709_ ), .A2(_01493_ ), .A3(_02566_ ), .ZN(_02567_ ) );
BUF_X2 _09801_ ( .A(_02362_ ), .Z(_02568_ ) );
NAND3_X1 _09802_ ( .A1(_01483_ ), .A2(\de_pc [4] ), .A3(_02568_ ), .ZN(_02569_ ) );
AND3_X1 _09803_ ( .A1(_02562_ ), .A2(_02567_ ), .A3(_02569_ ), .ZN(_02570_ ) );
OAI21_X1 _09804_ ( .A(_02561_ ), .B1(_02570_ ), .B2(_01570_ ), .ZN(_00149_ ) );
MUX2_X1 _09805_ ( .A(\u_exu.ecsr [3] ), .B(\ea_addr [3] ), .S(_01134_ ), .Z(_02571_ ) );
OAI22_X1 _09806_ ( .A1(_01730_ ), .A2(_01247_ ), .B1(_01144_ ), .B2(_02187_ ), .ZN(_02572_ ) );
AOI21_X1 _09807_ ( .A(_01237_ ), .B1(_01734_ ), .B2(_01735_ ), .ZN(_02573_ ) );
OR3_X2 _09808_ ( .A1(_02572_ ), .A2(_01524_ ), .A3(_02573_ ), .ZN(_02574_ ) );
AOI21_X1 _09809_ ( .A(_01254_ ), .B1(io_master_rready ), .B2(\io_master_rdata [3] ), .ZN(_02575_ ) );
INV_X1 _09810_ ( .A(\u_lsu.u_clint.mtime [35] ), .ZN(_02576_ ) );
INV_X4 _09811_ ( .A(\u_lsu.u_clint.mtime [3] ), .ZN(_02577_ ) );
MUX2_X1 _09812_ ( .A(_02576_ ), .B(_02577_ ), .S(_01733_ ), .Z(_02578_ ) );
OAI21_X1 _09813_ ( .A(_02575_ ), .B1(_01229_ ), .B2(_02578_ ), .ZN(_02579_ ) );
AND3_X2 _09814_ ( .A1(_02574_ ), .A2(_02430_ ), .A3(_02579_ ), .ZN(_02580_ ) );
MUX2_X2 _09815_ ( .A(_02571_ ), .B(_02580_ ), .S(fanout_net_10 ), .Z(\ar_data [3] ) );
AND2_X2 _09816_ ( .A1(\ar_data [3] ), .A2(_01311_ ), .ZN(_02581_ ) );
AOI22_X1 _09817_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01319_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02582_ ) );
AOI22_X1 _09818_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01330_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02583_ ) );
NAND3_X1 _09819_ ( .A1(_02582_ ), .A2(_01325_ ), .A3(_02583_ ), .ZN(_02584_ ) );
OAI211_X1 _09820_ ( .A(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01337_ ), .C1(_01871_ ), .C2(_01872_ ), .ZN(_02585_ ) );
INV_X1 _09821_ ( .A(\u_reg.rf[1][3] ), .ZN(_02586_ ) );
AOI21_X1 _09822_ ( .A(_01342_ ), .B1(_01344_ ), .B2(_02586_ ), .ZN(_02587_ ) );
NOR2_X1 _09823_ ( .A1(_01344_ ), .A2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02588_ ) );
OAI211_X1 _09824_ ( .A(_01026_ ), .B(_02585_ ), .C1(_02587_ ), .C2(_02588_ ), .ZN(_02589_ ) );
NAND3_X1 _09825_ ( .A1(_02584_ ), .A2(_01813_ ), .A3(_02589_ ), .ZN(_02590_ ) );
AOI22_X1 _09826_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01319_ ), .B1(_01321_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02591_ ) );
AOI22_X1 _09827_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01327_ ), .B1(_01330_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02592_ ) );
AOI21_X1 _09828_ ( .A(_01026_ ), .B1(_02591_ ), .B2(_02592_ ), .ZN(_02593_ ) );
AOI22_X1 _09829_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01319_ ), .B1(_01321_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02594_ ) );
AOI22_X1 _09830_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01327_ ), .B1(_01330_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02595_ ) );
AOI21_X1 _09831_ ( .A(_01325_ ), .B1(_02594_ ), .B2(_02595_ ), .ZN(_02596_ ) );
OAI21_X1 _09832_ ( .A(_01043_ ), .B1(_02593_ ), .B2(_02596_ ), .ZN(_02597_ ) );
AND3_X1 _09833_ ( .A1(_01312_ ), .A2(_02590_ ), .A3(_02597_ ), .ZN(_02598_ ) );
OAI21_X1 _09834_ ( .A(_01535_ ), .B1(_02581_ ), .B2(_02598_ ), .ZN(_02599_ ) );
OR2_X2 _09835_ ( .A1(_02599_ ), .A2(_01832_ ), .ZN(_02600_ ) );
AND4_X1 _09836_ ( .A1(\u_csr.csr[0][3] ), .A2(_01465_ ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_02601_ ) );
AOI21_X1 _09837_ ( .A(_02601_ ), .B1(_02494_ ), .B2(\u_csr.csr[1][3] ), .ZN(_02602_ ) );
INV_X1 _09838_ ( .A(_01641_ ), .ZN(_02603_ ) );
NAND4_X1 _09839_ ( .A1(_01651_ ), .A2(\u_csr.csr[2][3] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_02604_ ) );
OAI211_X1 _09840_ ( .A(_01591_ ), .B(\u_csr.csr[3][0] ), .C1(_00754_ ), .C2(_00857_ ), .ZN(_02605_ ) );
NOR3_X1 _09841_ ( .A1(_02605_ ), .A2(_01642_ ), .A3(_01643_ ), .ZN(_02606_ ) );
NOR2_X1 _09842_ ( .A1(_01645_ ), .A2(_02606_ ), .ZN(_02607_ ) );
NAND4_X1 _09843_ ( .A1(_02602_ ), .A2(_02603_ ), .A3(_02604_ ), .A4(_02607_ ), .ZN(_02608_ ) );
NAND2_X1 _09844_ ( .A1(_01575_ ), .A2(_02608_ ), .ZN(_02609_ ) );
NAND4_X1 _09845_ ( .A1(_01774_ ), .A2(_00830_ ), .A3(_00828_ ), .A4(_01715_ ), .ZN(_02610_ ) );
AOI21_X1 _09846_ ( .A(_01767_ ), .B1(_02609_ ), .B2(_02610_ ), .ZN(_02611_ ) );
AOI221_X4 _09847_ ( .A(_02611_ ), .B1(\de_pc [3] ), .B2(_01479_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_02612_ ) );
OR2_X1 _09848_ ( .A1(_02599_ ), .A2(_01483_ ), .ZN(_02613_ ) );
NOR2_X1 _09849_ ( .A1(_01496_ ), .A2(_00918_ ), .ZN(_02614_ ) );
AOI21_X1 _09850_ ( .A(_00888_ ), .B1(_00727_ ), .B2(_00895_ ), .ZN(_02615_ ) );
OR2_X1 _09851_ ( .A1(_02614_ ), .A2(_02615_ ), .ZN(_02616_ ) );
AOI221_X1 _09852_ ( .A(_01487_ ), .B1(\de_pc [3] ), .B2(_01491_ ), .C1(_01720_ ), .C2(_02616_ ), .ZN(_02617_ ) );
AOI221_X1 _09853_ ( .A(_02275_ ), .B1(_02600_ ), .B2(_02612_ ), .C1(_02613_ ), .C2(_02617_ ), .ZN(_00150_ ) );
MUX2_X1 _09854_ ( .A(\u_exu.ecsr [2] ), .B(\ea_addr [2] ), .S(_01134_ ), .Z(_02618_ ) );
AND3_X1 _09855_ ( .A1(_01798_ ), .A2(_01246_ ), .A3(_01800_ ), .ZN(_02619_ ) );
AOI21_X1 _09856_ ( .A(_02619_ ), .B1(_01236_ ), .B2(_01796_ ), .ZN(_02620_ ) );
NOR2_X1 _09857_ ( .A1(_02233_ ), .A2(_01144_ ), .ZN(_02621_ ) );
INV_X1 _09858_ ( .A(_02621_ ), .ZN(_02622_ ) );
AND3_X1 _09859_ ( .A1(_02620_ ), .A2(_01254_ ), .A3(_02622_ ), .ZN(_02623_ ) );
AND2_X1 _09860_ ( .A1(io_master_rready ), .A2(\io_master_rdata [2] ), .ZN(_02624_ ) );
AND3_X1 _09861_ ( .A1(_01212_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ), .A3(_01213_ ), .ZN(_02625_ ) );
INV_X1 _09862_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_28_A_$_ANDNOT__Y_B ), .ZN(_02626_ ) );
AOI21_X1 _09863_ ( .A(_02626_ ), .B1(_01669_ ), .B2(_01213_ ), .ZN(_02627_ ) );
NOR3_X1 _09864_ ( .A1(_02625_ ), .A2(_02627_ ), .A3(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ), .ZN(_02628_ ) );
AND2_X1 _09865_ ( .A1(_01526_ ), .A2(_02628_ ), .ZN(_02629_ ) );
NOR3_X1 _09866_ ( .A1(_02624_ ), .A2(_01254_ ), .A3(_02629_ ), .ZN(_02630_ ) );
NOR3_X1 _09867_ ( .A1(_02623_ ), .A2(_02365_ ), .A3(_02630_ ), .ZN(_02631_ ) );
MUX2_X1 _09868_ ( .A(_02618_ ), .B(_02631_ ), .S(fanout_net_10 ), .Z(\ar_data [2] ) );
NAND2_X1 _09869_ ( .A1(\ar_data [2] ), .A2(_01318_ ), .ZN(_02632_ ) );
AOI22_X1 _09870_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02633_ ) );
AOI22_X1 _09871_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02634_ ) );
AOI21_X1 _09872_ ( .A(_01633_ ), .B1(_02633_ ), .B2(_02634_ ), .ZN(_02635_ ) );
AOI22_X1 _09873_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02636_ ) );
AOI22_X1 _09874_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01752_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02637_ ) );
AOI21_X1 _09875_ ( .A(_01557_ ), .B1(_02636_ ), .B2(_02637_ ), .ZN(_02638_ ) );
OAI21_X1 _09876_ ( .A(_01366_ ), .B1(_02635_ ), .B2(_02638_ ), .ZN(_02639_ ) );
OAI211_X1 _09877_ ( .A(_01694_ ), .B(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C1(_01871_ ), .C2(_01872_ ), .ZN(_02640_ ) );
OAI211_X1 _09878_ ( .A(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(_02243_ ), .C1(_01871_ ), .C2(_01872_ ), .ZN(_02641_ ) );
NAND2_X1 _09879_ ( .A1(_02640_ ), .A2(_02641_ ), .ZN(_02642_ ) );
MUX2_X1 _09880_ ( .A(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_02243_ ), .Z(_02643_ ) );
AOI211_X1 _09881_ ( .A(_01354_ ), .B(_02642_ ), .C1(_02021_ ), .C2(_02643_ ), .ZN(_02644_ ) );
OAI21_X1 _09882_ ( .A(_02243_ ), .B1(_01545_ ), .B2(\u_reg.rf[1][2] ), .ZN(_02645_ ) );
OAI21_X1 _09883_ ( .A(_02645_ ), .B1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01551_ ), .ZN(_02646_ ) );
OAI211_X1 _09884_ ( .A(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01547_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_02647_ ) );
NAND3_X1 _09885_ ( .A1(_02646_ ), .A2(_01354_ ), .A3(_02647_ ), .ZN(_02648_ ) );
NAND2_X1 _09886_ ( .A1(_02648_ ), .A2(_01334_ ), .ZN(_02649_ ) );
OAI21_X1 _09887_ ( .A(_02639_ ), .B1(_02644_ ), .B2(_02649_ ), .ZN(_02650_ ) );
OR2_X1 _09888_ ( .A1(_01318_ ), .A2(_02650_ ), .ZN(_02651_ ) );
AOI21_X1 _09889_ ( .A(_01805_ ), .B1(_02632_ ), .B2(_02651_ ), .ZN(_02652_ ) );
AND2_X1 _09890_ ( .A1(_02652_ ), .A2(_01371_ ), .ZN(_02653_ ) );
NAND3_X1 _09891_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][2] ), .A3(_01455_ ), .ZN(_02654_ ) );
NAND4_X1 _09892_ ( .A1(_01582_ ), .A2(\u_csr.csr[2][2] ), .A3(_00754_ ), .A4(_01591_ ), .ZN(_02655_ ) );
AND2_X1 _09893_ ( .A1(_01457_ ), .A2(_01460_ ), .ZN(_02656_ ) );
AOI22_X1 _09894_ ( .A1(_02656_ ), .A2(\u_csr.csr[0][2] ), .B1(_01644_ ), .B2(_01587_ ), .ZN(_02657_ ) );
AND2_X1 _09895_ ( .A1(_02655_ ), .A2(_02657_ ), .ZN(_02658_ ) );
AOI21_X1 _09896_ ( .A(_02492_ ), .B1(_02654_ ), .B2(_02658_ ), .ZN(_02659_ ) );
AOI22_X1 _09897_ ( .A1(\u_idu.imm_auipc_lui [31] ), .A2(_01385_ ), .B1(_01434_ ), .B2(\u_idu.imm_auipc_lui [30] ), .ZN(_02660_ ) );
OAI22_X1 _09898_ ( .A1(_01399_ ), .A2(_00887_ ), .B1(_01391_ ), .B2(_00734_ ), .ZN(_02661_ ) );
AOI221_X4 _09899_ ( .A(_02661_ ), .B1(\u_idu.imm_auipc_lui [25] ), .B2(_01414_ ), .C1(_00881_ ), .C2(_01431_ ), .ZN(_02662_ ) );
AOI22_X1 _09900_ ( .A1(_02660_ ), .A2(_02662_ ), .B1(_00760_ ), .B2(ea_err ), .ZN(_02663_ ) );
AOI221_X4 _09901_ ( .A(_01395_ ), .B1(\u_idu.imm_auipc_lui [28] ), .B2(_01388_ ), .C1(_00656_ ), .C2(_01413_ ), .ZN(_02664_ ) );
AOI22_X1 _09902_ ( .A1(_01433_ ), .A2(_00861_ ), .B1(_01430_ ), .B2(\u_idu.imm_auipc_lui [29] ), .ZN(_02665_ ) );
AND4_X1 _09903_ ( .A1(_01436_ ), .A2(_02504_ ), .A3(_01393_ ), .A4(_01402_ ), .ZN(_02666_ ) );
NAND4_X1 _09904_ ( .A1(_01381_ ), .A2(_02664_ ), .A3(_02665_ ), .A4(_02666_ ), .ZN(_02667_ ) );
OAI22_X1 _09905_ ( .A1(_01410_ ), .A2(_00886_ ), .B1(\u_idu.imm_auipc_lui [28] ), .B2(_01388_ ), .ZN(_02668_ ) );
AOI211_X1 _09906_ ( .A(_02663_ ), .B(_02667_ ), .C1(_00640_ ), .C2(_02668_ ), .ZN(_02669_ ) );
INV_X1 _09907_ ( .A(_01397_ ), .ZN(_02670_ ) );
AND3_X1 _09908_ ( .A1(_02669_ ), .A2(_02505_ ), .A3(_02670_ ), .ZN(_02671_ ) );
AND3_X1 _09909_ ( .A1(_02671_ ), .A2(_01408_ ), .A3(_01383_ ), .ZN(_02672_ ) );
NAND3_X1 _09910_ ( .A1(_02672_ ), .A2(_01428_ ), .A3(_01379_ ), .ZN(_02673_ ) );
AOI211_X1 _09911_ ( .A(_01441_ ), .B(_02673_ ), .C1(_00831_ ), .C2(_00832_ ), .ZN(_02674_ ) );
NOR2_X1 _09912_ ( .A1(_02659_ ), .A2(_02674_ ), .ZN(_02675_ ) );
INV_X1 _09913_ ( .A(\de_pc [2] ), .ZN(_02676_ ) );
OAI22_X1 _09914_ ( .A1(_02675_ ), .A2(_01375_ ), .B1(_02676_ ), .B2(_01478_ ), .ZN(_02677_ ) );
OAI21_X1 _09915_ ( .A(_01855_ ), .B1(_02653_ ), .B2(_02677_ ), .ZN(_02678_ ) );
NAND2_X1 _09916_ ( .A1(_02652_ ), .A2(_01485_ ), .ZN(_02679_ ) );
AND2_X1 _09917_ ( .A1(_02563_ ), .A2(\u_idu.imm_branch [2] ), .ZN(_02680_ ) );
AOI21_X1 _09918_ ( .A(_00890_ ), .B1(_00727_ ), .B2(_00895_ ), .ZN(_02681_ ) );
NOR2_X1 _09919_ ( .A1(_02680_ ), .A2(_02681_ ), .ZN(_02682_ ) );
INV_X1 _09920_ ( .A(_02682_ ), .ZN(_02683_ ) );
NAND3_X1 _09921_ ( .A1(_00709_ ), .A2(_01493_ ), .A3(_02683_ ), .ZN(_02684_ ) );
NAND3_X1 _09922_ ( .A1(_01483_ ), .A2(\de_pc [2] ), .A3(_02362_ ), .ZN(_02685_ ) );
AND3_X1 _09923_ ( .A1(_02679_ ), .A2(_02684_ ), .A3(_02685_ ), .ZN(_02686_ ) );
OAI21_X1 _09924_ ( .A(_02678_ ), .B1(_02686_ ), .B2(_01570_ ), .ZN(_00151_ ) );
AOI22_X1 _09925_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01806_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02687_ ) );
AOI22_X1 _09926_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02688_ ) );
AOI21_X1 _09927_ ( .A(_01558_ ), .B1(_02687_ ), .B2(_02688_ ), .ZN(_02689_ ) );
AOI22_X1 _09928_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01537_ ), .B1(_01807_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02690_ ) );
AOI22_X1 _09929_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01541_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02691_ ) );
AOI21_X1 _09930_ ( .A(_01326_ ), .B1(_02690_ ), .B2(_02691_ ), .ZN(_02692_ ) );
OAI21_X1 _09931_ ( .A(_01822_ ), .B1(_02689_ ), .B2(_02692_ ), .ZN(_02693_ ) );
AOI22_X1 _09932_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02694_ ) );
AOI22_X1 _09933_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02695_ ) );
AND3_X1 _09934_ ( .A1(_02694_ ), .A2(_01756_ ), .A3(_02695_ ), .ZN(_02696_ ) );
OR2_X1 _09935_ ( .A1(_02696_ ), .A2(_01366_ ), .ZN(_02697_ ) );
OAI21_X1 _09936_ ( .A(_01338_ ), .B1(_01545_ ), .B2(\u_reg.rf[1][28] ), .ZN(_02698_ ) );
INV_X1 _09937_ ( .A(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02699_ ) );
OAI21_X1 _09938_ ( .A(_02699_ ), .B1(_01871_ ), .B2(_01872_ ), .ZN(_02700_ ) );
AOI221_X4 _09939_ ( .A(_01325_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(_02698_ ), .C2(_02700_ ), .ZN(_02701_ ) );
OAI21_X1 _09940_ ( .A(_02693_ ), .B1(_02697_ ), .B2(_02701_ ), .ZN(_02702_ ) );
AOI21_X1 _09941_ ( .A(_01805_ ), .B1(_01856_ ), .B2(_02702_ ), .ZN(_02703_ ) );
AND3_X1 _09942_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [28] ), .ZN(_02704_ ) );
AOI211_X1 _09943_ ( .A(fanout_net_10 ), .B(_02704_ ), .C1(\ea_addr [28] ), .C2(_01521_ ), .ZN(_02705_ ) );
AOI21_X4 _09944_ ( .A(_01523_ ), .B1(_01525_ ), .B2(_01675_ ), .ZN(_02706_ ) );
AOI21_X4 _09945_ ( .A(_02705_ ), .B1(_02706_ ), .B2(fanout_net_10 ), .ZN(\ar_data [28] ) );
OAI21_X2 _09946_ ( .A(_02703_ ), .B1(\ar_data [28] ), .B2(_01856_ ), .ZN(_02707_ ) );
NOR2_X1 _09947_ ( .A1(_02707_ ), .A2(_01833_ ), .ZN(_02708_ ) );
AND3_X1 _09948_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][28] ), .A3(_01462_ ), .ZN(_02709_ ) );
AOI21_X1 _09949_ ( .A(_02709_ ), .B1(_01584_ ), .B2(_01588_ ), .ZN(_02710_ ) );
NAND3_X1 _09950_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][28] ), .A3(_01579_ ), .ZN(_02711_ ) );
NAND4_X1 _09951_ ( .A1(_01579_ ), .A2(\u_csr.csr[2][28] ), .A3(_01653_ ), .A4(_01649_ ), .ZN(_02712_ ) );
NAND3_X1 _09952_ ( .A1(_02710_ ), .A2(_02711_ ), .A3(_02712_ ), .ZN(_02713_ ) );
NAND3_X1 _09953_ ( .A1(_01439_ ), .A2(_01597_ ), .A3(_02713_ ), .ZN(_02714_ ) );
NAND4_X1 _09954_ ( .A1(_01596_ ), .A2(_00838_ ), .A3(_00837_ ), .A4(_01597_ ), .ZN(_02715_ ) );
AND2_X1 _09955_ ( .A1(_02714_ ), .A2(_02715_ ), .ZN(_02716_ ) );
INV_X1 _09956_ ( .A(\de_pc [28] ), .ZN(_02717_ ) );
OAI22_X1 _09957_ ( .A1(_02716_ ), .A2(_01375_ ), .B1(_02717_ ), .B2(_01478_ ), .ZN(_02718_ ) );
OAI21_X1 _09958_ ( .A(_01855_ ), .B1(_02708_ ), .B2(_02718_ ), .ZN(_02719_ ) );
OAI22_X1 _09959_ ( .A1(_02707_ ), .A2(_01483_ ), .B1(_02717_ ), .B2(_01507_ ), .ZN(_02720_ ) );
NAND3_X1 _09960_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [28] ), .A3(_01512_ ), .ZN(_02721_ ) );
NAND3_X1 _09961_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_02721_ ), .ZN(_02722_ ) );
AOI21_X1 _09962_ ( .A(_02720_ ), .B1(_01495_ ), .B2(_02722_ ), .ZN(_02723_ ) );
OAI21_X1 _09963_ ( .A(_02719_ ), .B1(_02723_ ), .B2(_01570_ ), .ZN(_00152_ ) );
MUX2_X1 _09964_ ( .A(\u_exu.ecsr [1] ), .B(\ea_addr [1] ), .S(_01136_ ), .Z(_02724_ ) );
AOI21_X1 _09965_ ( .A(_01247_ ), .B1(_01881_ ), .B2(_01882_ ), .ZN(_02725_ ) );
AOI21_X1 _09966_ ( .A(_02725_ ), .B1(_02281_ ), .B2(_01236_ ), .ZN(_02726_ ) );
OAI21_X1 _09967_ ( .A(_01143_ ), .B1(_02276_ ), .B2(_02278_ ), .ZN(_02727_ ) );
NAND3_X1 _09968_ ( .A1(_02726_ ), .A2(_01277_ ), .A3(_02727_ ), .ZN(_02728_ ) );
OR2_X1 _09969_ ( .A1(_01733_ ), .A2(\u_lsu.u_clint.mtime [33] ), .ZN(_02729_ ) );
OAI211_X1 _09970_ ( .A(_01238_ ), .B(_02729_ ), .C1(\u_lsu.u_clint.mtime [1] ), .C2(_01249_ ), .ZN(_02730_ ) );
OAI21_X1 _09971_ ( .A(\io_master_rdata [1] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_02731_ ) );
NAND3_X1 _09972_ ( .A1(_02730_ ), .A2(_01524_ ), .A3(_02731_ ), .ZN(_02732_ ) );
AND3_X1 _09973_ ( .A1(_02728_ ), .A2(_02431_ ), .A3(_02732_ ), .ZN(_02733_ ) );
MUX2_X1 _09974_ ( .A(_02724_ ), .B(_02733_ ), .S(fanout_net_10 ), .Z(\ar_data [1] ) );
NAND2_X1 _09975_ ( .A1(\ar_data [1] ), .A2(_01318_ ), .ZN(_02734_ ) );
AND3_X1 _09976_ ( .A1(_01307_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01336_ ), .ZN(_02735_ ) );
AOI221_X4 _09977_ ( .A(_02735_ ), .B1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01540_ ), .C1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(_01757_ ), .ZN(_02736_ ) );
AOI21_X1 _09978_ ( .A(_01326_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02737_ ) );
AOI21_X1 _09979_ ( .A(_01334_ ), .B1(_02736_ ), .B2(_02737_ ), .ZN(_02738_ ) );
AOI22_X1 _09980_ ( .A1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_02012_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02739_ ) );
AOI22_X1 _09981_ ( .A1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02740_ ) );
NAND3_X1 _09982_ ( .A1(_02739_ ), .A2(_02015_ ), .A3(_02740_ ), .ZN(_02741_ ) );
NAND2_X1 _09983_ ( .A1(_02738_ ), .A2(_02741_ ), .ZN(_02742_ ) );
AOI22_X1 _09984_ ( .A1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_02012_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02743_ ) );
OAI211_X1 _09985_ ( .A(_01816_ ), .B(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_02744_ ) );
OAI211_X1 _09986_ ( .A(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(_01965_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_02745_ ) );
AND4_X1 _09987_ ( .A1(_02015_ ), .A2(_02743_ ), .A3(_02744_ ), .A4(_02745_ ), .ZN(_02746_ ) );
OAI211_X1 _09988_ ( .A(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01965_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_02747_ ) );
INV_X1 _09989_ ( .A(\u_reg.rf[1][1] ), .ZN(_02748_ ) );
AOI21_X1 _09990_ ( .A(_01816_ ), .B1(_02021_ ), .B2(_02748_ ), .ZN(_02749_ ) );
NOR2_X1 _09991_ ( .A1(_02021_ ), .A2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02750_ ) );
OAI211_X1 _09992_ ( .A(_01858_ ), .B(_02747_ ), .C1(_02749_ ), .C2(_02750_ ), .ZN(_02751_ ) );
NAND2_X1 _09993_ ( .A1(_02751_ ), .A2(_01814_ ), .ZN(_02752_ ) );
OAI211_X1 _09994_ ( .A(_01536_ ), .B(_02742_ ), .C1(_02746_ ), .C2(_02752_ ), .ZN(_02753_ ) );
AOI21_X1 _09995_ ( .A(_01805_ ), .B1(_02734_ ), .B2(_02753_ ), .ZN(_02754_ ) );
AND2_X1 _09996_ ( .A1(_02754_ ), .A2(_01371_ ), .ZN(_02755_ ) );
NAND4_X1 _09997_ ( .A1(_01584_ ), .A2(\u_csr.csr[2][1] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_02756_ ) );
INV_X1 _09998_ ( .A(_01645_ ), .ZN(_02757_ ) );
INV_X1 _09999_ ( .A(_02606_ ), .ZN(_02758_ ) );
NAND3_X1 _10000_ ( .A1(_02756_ ), .A2(_02757_ ), .A3(_02758_ ), .ZN(_02759_ ) );
NAND3_X1 _10001_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][1] ), .A3(_01579_ ), .ZN(_02760_ ) );
NAND3_X1 _10002_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][1] ), .A3(_01462_ ), .ZN(_02761_ ) );
NAND2_X1 _10003_ ( .A1(_02760_ ), .A2(_02761_ ), .ZN(_02762_ ) );
OAI21_X1 _10004_ ( .A(_01576_ ), .B1(_02759_ ), .B2(_02762_ ), .ZN(_02763_ ) );
AND4_X1 _10005_ ( .A1(_01379_ ), .A2(_02671_ ), .A3(_01408_ ), .A4(_01383_ ), .ZN(_02764_ ) );
NAND2_X1 _10006_ ( .A1(_00833_ ), .A2(_00834_ ), .ZN(_02765_ ) );
NAND4_X1 _10007_ ( .A1(_02764_ ), .A2(_02765_ ), .A3(_01597_ ), .A4(_01428_ ), .ZN(_02766_ ) );
AND2_X1 _10008_ ( .A1(_02763_ ), .A2(_02766_ ), .ZN(_02767_ ) );
INV_X1 _10009_ ( .A(\de_pc [1] ), .ZN(_02768_ ) );
OAI22_X1 _10010_ ( .A1(_02767_ ), .A2(_01375_ ), .B1(_02768_ ), .B2(_01478_ ), .ZN(_02769_ ) );
OAI21_X1 _10011_ ( .A(_01855_ ), .B1(_02755_ ), .B2(_02769_ ), .ZN(_02770_ ) );
NAND2_X1 _10012_ ( .A1(_02754_ ), .A2(_01485_ ), .ZN(_02771_ ) );
AND2_X1 _10013_ ( .A1(_02563_ ), .A2(\u_idu.imm_branch [1] ), .ZN(_02772_ ) );
CLKBUF_X2 _10014_ ( .A(_00978_ ), .Z(_02773_ ) );
BUF_X2 _10015_ ( .A(_02773_ ), .Z(_02774_ ) );
BUF_X2 _10016_ ( .A(_02774_ ), .Z(_02775_ ) );
BUF_X4 _10017_ ( .A(_02775_ ), .Z(_02776_ ) );
AOI21_X1 _10018_ ( .A(_02776_ ), .B1(_00727_ ), .B2(_00895_ ), .ZN(_02777_ ) );
NOR2_X1 _10019_ ( .A1(_02772_ ), .A2(_02777_ ), .ZN(_02778_ ) );
INV_X1 _10020_ ( .A(_02778_ ), .ZN(_02779_ ) );
NAND3_X1 _10021_ ( .A1(_00709_ ), .A2(_01493_ ), .A3(_02779_ ), .ZN(_02780_ ) );
NAND3_X1 _10022_ ( .A1(_01483_ ), .A2(\de_pc [1] ), .A3(_02362_ ), .ZN(_02781_ ) );
AND3_X1 _10023_ ( .A1(_02771_ ), .A2(_02780_ ), .A3(_02781_ ), .ZN(_02782_ ) );
OAI21_X1 _10024_ ( .A(_02770_ ), .B1(_02782_ ), .B2(_01570_ ), .ZN(_00153_ ) );
AOI22_X1 _10025_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01757_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02783_ ) );
AOI22_X1 _10026_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02784_ ) );
AOI21_X1 _10027_ ( .A(_00944_ ), .B1(_02783_ ), .B2(_02784_ ), .ZN(_02785_ ) );
OAI211_X1 _10028_ ( .A(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01338_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_02786_ ) );
INV_X1 _10029_ ( .A(\u_reg.rf[1][0] ), .ZN(_02787_ ) );
AOI21_X1 _10030_ ( .A(_01343_ ), .B1(_01551_ ), .B2(_02787_ ), .ZN(_02788_ ) );
NOR2_X1 _10031_ ( .A1(_01551_ ), .A2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02789_ ) );
OAI21_X1 _10032_ ( .A(_02786_ ), .B1(_02788_ ), .B2(_02789_ ), .ZN(_02790_ ) );
AOI211_X1 _10033_ ( .A(_01809_ ), .B(_02785_ ), .C1(_01334_ ), .C2(_02790_ ), .ZN(_02791_ ) );
AOI22_X1 _10034_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01320_ ), .B1(_01538_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02792_ ) );
AOI22_X1 _10035_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01559_ ), .B1(_01331_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02793_ ) );
AOI21_X1 _10036_ ( .A(_01813_ ), .B1(_02792_ ), .B2(_02793_ ), .ZN(_02794_ ) );
AOI22_X1 _10037_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02795_ ) );
AOI22_X1 _10038_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02796_ ) );
AOI21_X1 _10039_ ( .A(_01043_ ), .B1(_02795_ ), .B2(_02796_ ), .ZN(_02797_ ) );
NOR3_X1 _10040_ ( .A1(_02794_ ), .A2(_02797_ ), .A3(_01858_ ), .ZN(_02798_ ) );
OAI21_X1 _10041_ ( .A(_01313_ ), .B1(_02791_ ), .B2(_02798_ ), .ZN(_02799_ ) );
NAND4_X1 _10042_ ( .A1(_01239_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D [0] ), .A3(\io_master_araddr [3] ), .A4(_01524_ ), .ZN(_02800_ ) );
INV_X1 _10043_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A ), .ZN(_02801_ ) );
OAI211_X1 _10044_ ( .A(_01238_ ), .B(_02800_ ), .C1(_02801_ ), .C2(_01733_ ), .ZN(_02802_ ) );
OAI21_X1 _10045_ ( .A(\io_master_rdata [0] ), .B1(_01607_ ), .B2(_01608_ ), .ZN(_02803_ ) );
AOI21_X1 _10046_ ( .A(_01276_ ), .B1(_02802_ ), .B2(_02803_ ), .ZN(_02804_ ) );
NAND3_X1 _10047_ ( .A1(_01914_ ), .A2(_02004_ ), .A3(_01918_ ), .ZN(_02805_ ) );
NAND3_X1 _10048_ ( .A1(_01908_ ), .A2(_01236_ ), .A3(_01911_ ), .ZN(_02806_ ) );
OAI211_X1 _10049_ ( .A(_02805_ ), .B(_02806_ ), .C1(_01144_ ), .C2(_02324_ ), .ZN(_02807_ ) );
OAI21_X1 _10050_ ( .A(_02431_ ), .B1(_02804_ ), .B2(_02807_ ), .ZN(_02808_ ) );
NAND2_X1 _10051_ ( .A1(_02808_ ), .A2(fanout_net_10 ), .ZN(_02809_ ) );
MUX2_X1 _10052_ ( .A(\u_exu.ecsr [0] ), .B(\ea_addr [0] ), .S(_01134_ ), .Z(_02810_ ) );
OR2_X1 _10053_ ( .A1(_02810_ ), .A2(fanout_net_10 ), .ZN(_02811_ ) );
NAND4_X1 _10054_ ( .A1(_02809_ ), .A2(_01286_ ), .A3(_01310_ ), .A4(_02811_ ), .ZN(_02812_ ) );
AOI21_X1 _10055_ ( .A(_01317_ ), .B1(_02799_ ), .B2(_02812_ ), .ZN(_02813_ ) );
NAND2_X1 _10056_ ( .A1(_02813_ ), .A2(_01370_ ), .ZN(_02814_ ) );
AND4_X1 _10057_ ( .A1(\u_csr.csr[2][0] ), .A2(_01453_ ), .A3(_01465_ ), .A4(_01467_ ), .ZN(_02815_ ) );
NAND4_X1 _10058_ ( .A1(_01465_ ), .A2(\u_csr.csr[0][0] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_02816_ ) );
NAND3_X1 _10059_ ( .A1(_02757_ ), .A2(_02758_ ), .A3(_02816_ ), .ZN(_02817_ ) );
AOI211_X1 _10060_ ( .A(_02815_ ), .B(_02817_ ), .C1(\u_csr.csr[1][0] ), .C2(_02494_ ), .ZN(_02818_ ) );
NOR2_X1 _10061_ ( .A1(_02818_ ), .A2(_02492_ ), .ZN(_02819_ ) );
NAND2_X1 _10062_ ( .A1(_00835_ ), .A2(_00836_ ), .ZN(_02820_ ) );
AND3_X1 _10063_ ( .A1(_01472_ ), .A2(_02820_ ), .A3(_01442_ ), .ZN(_02821_ ) );
NOR2_X4 _10064_ ( .A1(_02819_ ), .A2(_02821_ ), .ZN(_02822_ ) );
NOR2_X1 _10065_ ( .A1(_02822_ ), .A2(_01375_ ), .ZN(_02823_ ) );
AOI221_X4 _10066_ ( .A(_02823_ ), .B1(\de_pc [0] ), .B2(_01479_ ), .C1(_01109_ ), .C2(_01105_ ), .ZN(_02824_ ) );
NAND2_X1 _10067_ ( .A1(_02813_ ), .A2(_01484_ ), .ZN(_02825_ ) );
NAND4_X1 _10068_ ( .A1(_00718_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(_00713_ ), .A4(_00683_ ), .ZN(_02826_ ) );
OAI21_X1 _10069_ ( .A(_02826_ ), .B1(_00898_ ), .B2(\u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ), .ZN(_02827_ ) );
AND3_X1 _10070_ ( .A1(_00691_ ), .A2(\u_idu.imm_branch [11] ), .A3(\u_idu.inst [5] ), .ZN(_02828_ ) );
AND3_X1 _10071_ ( .A1(_00672_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(_00677_ ), .ZN(_02829_ ) );
OR3_X1 _10072_ ( .A1(_02827_ ), .A2(_02828_ ), .A3(_02829_ ), .ZN(_02830_ ) );
AOI221_X4 _10073_ ( .A(_01056_ ), .B1(\de_pc [0] ), .B2(_01491_ ), .C1(_01720_ ), .C2(_02830_ ), .ZN(_02831_ ) );
AOI221_X1 _10074_ ( .A(_02275_ ), .B1(_02814_ ), .B2(_02824_ ), .C1(_02825_ ), .C2(_02831_ ), .ZN(_00154_ ) );
AND3_X1 _10075_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [27] ), .ZN(_02832_ ) );
AOI211_X1 _10076_ ( .A(fanout_net_10 ), .B(_02832_ ), .C1(\ea_addr [27] ), .C2(_01521_ ), .ZN(_02833_ ) );
AOI21_X4 _10077_ ( .A(_01523_ ), .B1(_01525_ ), .B2(_01736_ ), .ZN(_02834_ ) );
AOI21_X4 _10078_ ( .A(_02833_ ), .B1(_02834_ ), .B2(fanout_net_10 ), .ZN(\ar_data [27] ) );
NOR2_X2 _10079_ ( .A1(\ar_data [27] ), .A2(_01686_ ), .ZN(_02835_ ) );
AOI22_X1 _10080_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01017_ ), .B1(_01321_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02836_ ) );
AOI22_X1 _10081_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01327_ ), .B1(_01329_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02837_ ) );
AND3_X1 _10082_ ( .A1(_02836_ ), .A2(_01324_ ), .A3(_02837_ ), .ZN(_02838_ ) );
OAI21_X1 _10083_ ( .A(_01336_ ), .B1(_01292_ ), .B2(\u_reg.rf[1][27] ), .ZN(_02839_ ) );
INV_X1 _10084_ ( .A(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02840_ ) );
OAI21_X1 _10085_ ( .A(_02840_ ), .B1(_00933_ ), .B2(_00934_ ), .ZN(_02841_ ) );
AOI221_X4 _10086_ ( .A(_00948_ ), .B1(_01329_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(_02839_ ), .C2(_02841_ ), .ZN(_02842_ ) );
OR3_X1 _10087_ ( .A1(_02838_ ), .A2(_01043_ ), .A3(_02842_ ), .ZN(_02843_ ) );
AOI22_X1 _10088_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02844_ ) );
AOI22_X1 _10089_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02845_ ) );
NAND3_X1 _10090_ ( .A1(_02844_ ), .A2(_01335_ ), .A3(_02845_ ), .ZN(_02846_ ) );
AOI22_X1 _10091_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02847_ ) );
AOI22_X1 _10092_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02848_ ) );
NAND3_X1 _10093_ ( .A1(_02847_ ), .A2(_01633_ ), .A3(_02848_ ), .ZN(_02849_ ) );
NAND3_X1 _10094_ ( .A1(_02846_ ), .A2(_02849_ ), .A3(_01705_ ), .ZN(_02850_ ) );
AOI21_X1 _10095_ ( .A(_01688_ ), .B1(_02843_ ), .B2(_02850_ ), .ZN(_02851_ ) );
NOR3_X2 _10096_ ( .A1(_02835_ ), .A2(_01316_ ), .A3(_02851_ ), .ZN(_02852_ ) );
NAND2_X1 _10097_ ( .A1(_02852_ ), .A2(_01370_ ), .ZN(_02853_ ) );
AND3_X1 _10098_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][27] ), .A3(_01647_ ), .ZN(_02854_ ) );
AND3_X1 _10099_ ( .A1(_01457_ ), .A2(\u_csr.csr[0][27] ), .A3(_01460_ ), .ZN(_02855_ ) );
AOI21_X1 _10100_ ( .A(_02855_ ), .B1(_01583_ ), .B2(_01587_ ), .ZN(_02856_ ) );
NAND4_X1 _10101_ ( .A1(_01582_ ), .A2(\u_csr.csr[2][27] ), .A3(_00754_ ), .A4(_01591_ ), .ZN(_02857_ ) );
NAND2_X1 _10102_ ( .A1(_02856_ ), .A2(_02857_ ), .ZN(_02858_ ) );
OAI21_X1 _10103_ ( .A(_01575_ ), .B1(_02854_ ), .B2(_02858_ ), .ZN(_02859_ ) );
NAND4_X1 _10104_ ( .A1(_01774_ ), .A2(_00840_ ), .A3(_00839_ ), .A4(_01443_ ), .ZN(_02860_ ) );
AOI21_X1 _10105_ ( .A(_01767_ ), .B1(_02859_ ), .B2(_02860_ ), .ZN(_02861_ ) );
AOI221_X4 _10106_ ( .A(_02861_ ), .B1(\de_pc [27] ), .B2(_01479_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_02862_ ) );
NAND2_X1 _10107_ ( .A1(_02852_ ), .A2(_01484_ ), .ZN(_02863_ ) );
NAND3_X1 _10108_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [27] ), .A3(_01512_ ), .ZN(_02864_ ) );
AND3_X1 _10109_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_02864_ ), .ZN(_02865_ ) );
NOR2_X1 _10110_ ( .A1(_01509_ ), .A2(_02865_ ), .ZN(_02866_ ) );
AOI211_X1 _10111_ ( .A(_02866_ ), .B(_01057_ ), .C1(\de_pc [27] ), .C2(_01492_ ), .ZN(_02867_ ) );
AOI221_X1 _10112_ ( .A(_02275_ ), .B1(_02853_ ), .B2(_02862_ ), .C1(_02863_ ), .C2(_02867_ ), .ZN(_00155_ ) );
NAND3_X1 _10113_ ( .A1(_01545_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_01694_ ), .ZN(_02868_ ) );
NAND3_X1 _10114_ ( .A1(_01928_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_02243_ ), .ZN(_02869_ ) );
NAND2_X1 _10115_ ( .A1(_02868_ ), .A2(_02869_ ), .ZN(_02870_ ) );
NAND3_X1 _10116_ ( .A1(_01545_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_02243_ ), .ZN(_02871_ ) );
NAND2_X1 _10117_ ( .A1(_02871_ ), .A2(_01756_ ), .ZN(_02872_ ) );
AOI211_X1 _10118_ ( .A(_02870_ ), .B(_02872_ ), .C1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_02012_ ), .ZN(_02873_ ) );
OR2_X1 _10119_ ( .A1(_02873_ ), .A2(_01814_ ), .ZN(_02874_ ) );
AOI22_X1 _10120_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_02012_ ), .B1(_02013_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02875_ ) );
AOI22_X1 _10121_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_02016_ ), .B1(_02017_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02876_ ) );
AND3_X1 _10122_ ( .A1(_02875_ ), .A2(_01858_ ), .A3(_02876_ ), .ZN(_02877_ ) );
OAI21_X1 _10123_ ( .A(_01547_ ), .B1(_01546_ ), .B2(\u_reg.rf[1][26] ), .ZN(_02878_ ) );
OR2_X1 _10124_ ( .A1(_01928_ ), .A2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02879_ ) );
AOI221_X4 _10125_ ( .A(_01756_ ), .B1(_01810_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C1(_02878_ ), .C2(_02879_ ), .ZN(_02880_ ) );
AOI22_X1 _10126_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01750_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02881_ ) );
AOI22_X1 _10127_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01752_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02882_ ) );
AND3_X1 _10128_ ( .A1(_02881_ ), .A2(_01756_ ), .A3(_02882_ ), .ZN(_02883_ ) );
OR2_X1 _10129_ ( .A1(_02883_ ), .A2(_01822_ ), .ZN(_02884_ ) );
OAI22_X1 _10130_ ( .A1(_02874_ ), .A2(_02877_ ), .B1(_02880_ ), .B2(_02884_ ), .ZN(_02885_ ) );
AOI21_X1 _10131_ ( .A(_01805_ ), .B1(_01856_ ), .B2(_02885_ ), .ZN(_02886_ ) );
AND3_X1 _10132_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [26] ), .ZN(_02887_ ) );
AOI211_X1 _10133_ ( .A(fanout_net_10 ), .B(_02887_ ), .C1(\ea_addr [26] ), .C2(_01521_ ), .ZN(_02888_ ) );
AOI21_X4 _10134_ ( .A(_01523_ ), .B1(_01525_ ), .B2(_01796_ ), .ZN(_02889_ ) );
AOI21_X4 _10135_ ( .A(_02888_ ), .B1(_02889_ ), .B2(fanout_net_10 ), .ZN(\ar_data [26] ) );
OAI21_X1 _10136_ ( .A(_02886_ ), .B1(\ar_data [26] ), .B2(_01856_ ), .ZN(_02890_ ) );
NOR2_X1 _10137_ ( .A1(_02890_ ), .A2(_01833_ ), .ZN(_02891_ ) );
NAND3_X1 _10138_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][26] ), .A3(_01579_ ), .ZN(_02892_ ) );
NAND4_X1 _10139_ ( .A1(_01584_ ), .A2(\u_csr.csr[2][26] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_02893_ ) );
NAND3_X1 _10140_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][26] ), .A3(_01462_ ), .ZN(_02894_ ) );
AND2_X1 _10141_ ( .A1(_02893_ ), .A2(_02894_ ), .ZN(_02895_ ) );
AOI21_X1 _10142_ ( .A(_02492_ ), .B1(_02892_ ), .B2(_02895_ ), .ZN(_02896_ ) );
AOI211_X1 _10143_ ( .A(_01441_ ), .B(_02673_ ), .C1(_00841_ ), .C2(_00842_ ), .ZN(_02897_ ) );
NOR2_X1 _10144_ ( .A1(_02896_ ), .A2(_02897_ ), .ZN(_02898_ ) );
INV_X1 _10145_ ( .A(\de_pc [26] ), .ZN(_02899_ ) );
OAI22_X1 _10146_ ( .A1(_02898_ ), .A2(_01843_ ), .B1(_02899_ ), .B2(_01845_ ), .ZN(_02900_ ) );
OAI21_X1 _10147_ ( .A(_01070_ ), .B1(_02891_ ), .B2(_02900_ ), .ZN(_02901_ ) );
BUF_X2 _10148_ ( .A(_01569_ ), .Z(_00302_ ) );
NOR2_X1 _10149_ ( .A1(_02890_ ), .A2(_01848_ ), .ZN(_02902_ ) );
NAND3_X1 _10150_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [26] ), .A3(_01512_ ), .ZN(_02903_ ) );
AND3_X1 _10151_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_02903_ ), .ZN(_02904_ ) );
OAI22_X1 _10152_ ( .A1(_01849_ ), .A2(_02899_ ), .B1(_01509_ ), .B2(_02904_ ), .ZN(_02905_ ) );
OAI21_X1 _10153_ ( .A(_00302_ ), .B1(_02902_ ), .B2(_02905_ ), .ZN(_02906_ ) );
NAND2_X1 _10154_ ( .A1(_02901_ ), .A2(_02906_ ), .ZN(_00156_ ) );
AND3_X1 _10155_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [25] ), .ZN(_02907_ ) );
AOI211_X1 _10156_ ( .A(fanout_net_10 ), .B(_02907_ ), .C1(\ea_addr [25] ), .C2(_01136_ ), .ZN(_02908_ ) );
AOI21_X4 _10157_ ( .A(_01523_ ), .B1(_01525_ ), .B2(_02281_ ), .ZN(_02909_ ) );
AOI21_X4 _10158_ ( .A(_02908_ ), .B1(_02909_ ), .B2(fanout_net_10 ), .ZN(\ar_data [25] ) );
NOR2_X2 _10159_ ( .A1(\ar_data [25] ), .A2(_01686_ ), .ZN(_02910_ ) );
AOI22_X1 _10160_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01351_ ), .B1(_01352_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02911_ ) );
AOI22_X1 _10161_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01328_ ), .B1(_01355_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02912_ ) );
NAND3_X1 _10162_ ( .A1(_02911_ ), .A2(_01361_ ), .A3(_02912_ ), .ZN(_02913_ ) );
NAND3_X1 _10163_ ( .A1(_01546_ ), .A2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01547_ ), .ZN(_02914_ ) );
OR3_X1 _10164_ ( .A1(_01871_ ), .A2(\u_reg.rf[1][25] ), .A3(_01872_ ), .ZN(_02915_ ) );
OAI21_X1 _10165_ ( .A(_01343_ ), .B1(_01345_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02916_ ) );
NAND4_X1 _10166_ ( .A1(_02914_ ), .A2(_01335_ ), .A3(_02915_ ), .A4(_02916_ ), .ZN(_02917_ ) );
NAND3_X1 _10167_ ( .A1(_02913_ ), .A2(_01813_ ), .A3(_02917_ ), .ZN(_02918_ ) );
AOI22_X1 _10168_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01358_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02919_ ) );
AOI22_X1 _10169_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01362_ ), .B1(_01363_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02920_ ) );
NAND3_X1 _10170_ ( .A1(_02919_ ), .A2(_01335_ ), .A3(_02920_ ), .ZN(_02921_ ) );
AOI22_X1 _10171_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01749_ ), .B1(_01359_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02922_ ) );
AOI22_X1 _10172_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01634_ ), .B1(_01753_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02923_ ) );
NAND3_X1 _10173_ ( .A1(_02922_ ), .A2(_01633_ ), .A3(_02923_ ), .ZN(_02924_ ) );
NAND3_X1 _10174_ ( .A1(_02921_ ), .A2(_02924_ ), .A3(_01705_ ), .ZN(_02925_ ) );
AOI21_X1 _10175_ ( .A(_01688_ ), .B1(_02918_ ), .B2(_02925_ ), .ZN(_02926_ ) );
NOR3_X2 _10176_ ( .A1(_02910_ ), .A2(_01316_ ), .A3(_02926_ ), .ZN(_02927_ ) );
NAND2_X1 _10177_ ( .A1(_02927_ ), .A2(_01370_ ), .ZN(_02928_ ) );
AND3_X1 _10178_ ( .A1(_01451_ ), .A2(\u_csr.csr[1][25] ), .A3(_01647_ ), .ZN(_02929_ ) );
NAND4_X1 _10179_ ( .A1(_01582_ ), .A2(\u_csr.csr[2][25] ), .A3(_00754_ ), .A4(_01591_ ), .ZN(_02930_ ) );
NAND3_X1 _10180_ ( .A1(_01458_ ), .A2(\u_csr.csr[0][25] ), .A3(_01461_ ), .ZN(_02931_ ) );
NAND2_X1 _10181_ ( .A1(_02930_ ), .A2(_02931_ ), .ZN(_02932_ ) );
OAI21_X1 _10182_ ( .A(_01575_ ), .B1(_02929_ ), .B2(_02932_ ), .ZN(_02933_ ) );
NAND4_X1 _10183_ ( .A1(_01774_ ), .A2(_00844_ ), .A3(_00843_ ), .A4(_01443_ ), .ZN(_02934_ ) );
AOI21_X1 _10184_ ( .A(_01767_ ), .B1(_02933_ ), .B2(_02934_ ), .ZN(_02935_ ) );
AOI221_X4 _10185_ ( .A(_02935_ ), .B1(\de_pc [25] ), .B2(_01479_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_02936_ ) );
NAND2_X1 _10186_ ( .A1(_02927_ ), .A2(_01484_ ), .ZN(_02937_ ) );
NAND3_X1 _10187_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [25] ), .A3(_01512_ ), .ZN(_02938_ ) );
NAND3_X1 _10188_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_02938_ ), .ZN(_02939_ ) );
AOI221_X1 _10189_ ( .A(_01056_ ), .B1(\de_pc [25] ), .B2(_01491_ ), .C1(_01720_ ), .C2(_02939_ ), .ZN(_02940_ ) );
AOI221_X1 _10190_ ( .A(_02275_ ), .B1(_02928_ ), .B2(_02936_ ), .C1(_02937_ ), .C2(_02940_ ), .ZN(_00157_ ) );
MUX2_X1 _10191_ ( .A(\u_exu.ecsr [24] ), .B(\ea_addr [24] ), .S(_01135_ ), .Z(_02941_ ) );
NOR2_X1 _10192_ ( .A1(_02941_ ), .A2(fanout_net_10 ), .ZN(_02942_ ) );
AOI21_X4 _10193_ ( .A(_01523_ ), .B1(_01525_ ), .B2(_01912_ ), .ZN(_02943_ ) );
AOI21_X2 _10194_ ( .A(_02942_ ), .B1(_02943_ ), .B2(fanout_net_10 ), .ZN(\ar_data [24] ) );
OR2_X2 _10195_ ( .A1(\ar_data [24] ), .A2(_01313_ ), .ZN(_02944_ ) );
NAND3_X1 _10196_ ( .A1(_01307_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01336_ ), .ZN(_02945_ ) );
INV_X1 _10197_ ( .A(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02946_ ) );
INV_X1 _10198_ ( .A(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02947_ ) );
OAI221_X1 _10199_ ( .A(_02945_ ), .B1(_02408_ ), .B2(_02946_ ), .C1(_02403_ ), .C2(_02947_ ), .ZN(_02948_ ) );
AND3_X1 _10200_ ( .A1(_01292_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_01342_ ), .ZN(_02949_ ) );
OR3_X1 _10201_ ( .A1(_02948_ ), .A2(_01026_ ), .A3(_02949_ ), .ZN(_02950_ ) );
AOI22_X1 _10202_ ( .A1(_01352_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01752_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02951_ ) );
NAND3_X1 _10203_ ( .A1(_01345_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01343_ ), .ZN(_02952_ ) );
NAND3_X1 _10204_ ( .A1(_01546_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01338_ ), .ZN(_02953_ ) );
NAND3_X1 _10205_ ( .A1(_02951_ ), .A2(_02952_ ), .A3(_02953_ ), .ZN(_02954_ ) );
OAI211_X1 _10206_ ( .A(_02950_ ), .B(_01366_ ), .C1(_01809_ ), .C2(_02954_ ), .ZN(_02955_ ) );
OAI211_X1 _10207_ ( .A(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01547_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_02956_ ) );
AOI21_X1 _10208_ ( .A(_01551_ ), .B1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01816_ ), .ZN(_02957_ ) );
INV_X1 _10209_ ( .A(\u_reg.rf[1][24] ), .ZN(_02958_ ) );
AOI21_X1 _10210_ ( .A(_02958_ ), .B1(_00936_ ), .B2(_00937_ ), .ZN(_02959_ ) );
OAI21_X1 _10211_ ( .A(_02956_ ), .B1(_02957_ ), .B2(_02959_ ), .ZN(_02960_ ) );
NOR2_X1 _10212_ ( .A1(_02960_ ), .A2(_02015_ ), .ZN(_02961_ ) );
NAND3_X1 _10213_ ( .A1(_01292_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_01342_ ), .ZN(_02962_ ) );
NAND3_X1 _10214_ ( .A1(_01307_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01336_ ), .ZN(_02963_ ) );
NAND2_X1 _10215_ ( .A1(_02962_ ), .A2(_02963_ ), .ZN(_02964_ ) );
NAND3_X1 _10216_ ( .A1(_01292_ ), .A2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01336_ ), .ZN(_02965_ ) );
NAND2_X1 _10217_ ( .A1(_02965_ ), .A2(_01324_ ), .ZN(_02966_ ) );
AOI211_X1 _10218_ ( .A(_02964_ ), .B(_02966_ ), .C1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_01757_ ), .ZN(_02967_ ) );
AOI21_X1 _10219_ ( .A(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_B ), .B1(_00932_ ), .B2(_00705_ ), .ZN(_02968_ ) );
OR3_X1 _10220_ ( .A1(_02967_ ), .A2(_00747_ ), .A3(_02968_ ), .ZN(_02969_ ) );
OAI21_X1 _10221_ ( .A(_02955_ ), .B1(_02961_ ), .B2(_02969_ ), .ZN(_02970_ ) );
AOI21_X1 _10222_ ( .A(_01316_ ), .B1(_01536_ ), .B2(_02970_ ), .ZN(_02971_ ) );
NAND3_X1 _10223_ ( .A1(_02944_ ), .A2(_01370_ ), .A3(_02971_ ), .ZN(_02972_ ) );
NAND4_X1 _10224_ ( .A1(_01651_ ), .A2(\u_csr.csr[2][24] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_02973_ ) );
NAND3_X1 _10225_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][24] ), .A3(_01651_ ), .ZN(_02974_ ) );
NAND4_X1 _10226_ ( .A1(_01653_ ), .A2(\u_csr.csr[0][24] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_02975_ ) );
NAND4_X1 _10227_ ( .A1(_01646_ ), .A2(_02973_ ), .A3(_02974_ ), .A4(_02975_ ), .ZN(_02976_ ) );
NAND2_X1 _10228_ ( .A1(_01575_ ), .A2(_02976_ ), .ZN(_02977_ ) );
NAND4_X1 _10229_ ( .A1(_01472_ ), .A2(_00846_ ), .A3(_00845_ ), .A4(_01443_ ), .ZN(_02978_ ) );
AOI21_X1 _10230_ ( .A(_01374_ ), .B1(_02977_ ), .B2(_02978_ ), .ZN(_02979_ ) );
AOI221_X4 _10231_ ( .A(_02979_ ), .B1(\de_pc [24] ), .B2(_01479_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_02980_ ) );
NAND3_X1 _10232_ ( .A1(_02944_ ), .A2(_01484_ ), .A3(_02971_ ), .ZN(_02981_ ) );
NAND3_X1 _10233_ ( .A1(_00713_ ), .A2(\u_idu.imm_auipc_lui [24] ), .A3(_00714_ ), .ZN(_02982_ ) );
AND3_X1 _10234_ ( .A1(_01498_ ), .A2(_01516_ ), .A3(_02982_ ), .ZN(_02983_ ) );
NOR2_X1 _10235_ ( .A1(_01509_ ), .A2(_02983_ ), .ZN(_02984_ ) );
AOI211_X1 _10236_ ( .A(_02984_ ), .B(_01057_ ), .C1(\de_pc [24] ), .C2(_01492_ ), .ZN(_02985_ ) );
AOI221_X1 _10237_ ( .A(_02275_ ), .B1(_02972_ ), .B2(_02980_ ), .C1(_02981_ ), .C2(_02985_ ), .ZN(_00158_ ) );
NAND3_X1 _10238_ ( .A1(_01545_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_01694_ ), .ZN(_02986_ ) );
NAND3_X1 _10239_ ( .A1(_01344_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01337_ ), .ZN(_02987_ ) );
NAND2_X1 _10240_ ( .A1(_02986_ ), .A2(_02987_ ), .ZN(_02988_ ) );
NAND3_X1 _10241_ ( .A1(_01545_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01337_ ), .ZN(_02989_ ) );
NAND2_X1 _10242_ ( .A1(_02989_ ), .A2(_01325_ ), .ZN(_02990_ ) );
AOI211_X1 _10243_ ( .A(_02988_ ), .B(_02990_ ), .C1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_02012_ ), .ZN(_02991_ ) );
AOI22_X1 _10244_ ( .A1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01319_ ), .B1(_01758_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02992_ ) );
AOI22_X1 _10245_ ( .A1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_01540_ ), .B1(_01760_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02993_ ) );
AND3_X1 _10246_ ( .A1(_02992_ ), .A2(_01557_ ), .A3(_02993_ ), .ZN(_02994_ ) );
OR3_X1 _10247_ ( .A1(_02991_ ), .A2(_01334_ ), .A3(_02994_ ), .ZN(_02995_ ) );
NAND3_X1 _10248_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_01816_ ), .ZN(_02996_ ) );
NAND3_X1 _10249_ ( .A1(_02021_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01965_ ), .ZN(_02997_ ) );
NAND2_X1 _10250_ ( .A1(_02996_ ), .A2(_02997_ ), .ZN(_02998_ ) );
NAND3_X1 _10251_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01965_ ), .ZN(_02999_ ) );
NAND2_X1 _10252_ ( .A1(_02999_ ), .A2(_01809_ ), .ZN(_03000_ ) );
AOI211_X1 _10253_ ( .A(_02998_ ), .B(_03000_ ), .C1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_02012_ ), .ZN(_03001_ ) );
OAI211_X1 _10254_ ( .A(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(_01965_ ), .C1(_01339_ ), .C2(_01340_ ), .ZN(_03002_ ) );
INV_X1 _10255_ ( .A(\u_reg.rf[1][23] ), .ZN(_03003_ ) );
AOI21_X1 _10256_ ( .A(_01816_ ), .B1(_02021_ ), .B2(_03003_ ), .ZN(_03004_ ) );
NOR2_X1 _10257_ ( .A1(_02021_ ), .A2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03005_ ) );
OAI21_X1 _10258_ ( .A(_03002_ ), .B1(_03004_ ), .B2(_03005_ ), .ZN(_03006_ ) );
OAI21_X1 _10259_ ( .A(_01814_ ), .B1(_03006_ ), .B2(_02015_ ), .ZN(_03007_ ) );
OAI21_X1 _10260_ ( .A(_02995_ ), .B1(_03001_ ), .B2(_03007_ ), .ZN(_03008_ ) );
AOI21_X1 _10261_ ( .A(_01805_ ), .B1(_01856_ ), .B2(_03008_ ), .ZN(_03009_ ) );
AND3_X1 _10262_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [23] ), .ZN(_03010_ ) );
AOI211_X1 _10263_ ( .A(fanout_net_10 ), .B(_03010_ ), .C1(\ea_addr [23] ), .C2(_01521_ ), .ZN(_03011_ ) );
NAND3_X1 _10264_ ( .A1(_01250_ ), .A2(_01524_ ), .A3(_01251_ ), .ZN(_03012_ ) );
AND3_X1 _10265_ ( .A1(_01243_ ), .A2(\io_master_araddr [0] ), .A3(_01244_ ), .ZN(_03013_ ) );
NOR4_X1 _10266_ ( .A1(_03013_ ), .A2(\io_master_araddr [1] ), .A3(_01274_ ), .A4(_01275_ ), .ZN(_03014_ ) );
AOI21_X4 _10267_ ( .A(_01523_ ), .B1(_03012_ ), .B2(_03014_ ), .ZN(_03015_ ) );
AOI21_X4 _10268_ ( .A(_03011_ ), .B1(_03015_ ), .B2(fanout_net_10 ), .ZN(\ar_data [23] ) );
OAI21_X1 _10269_ ( .A(_03009_ ), .B1(\ar_data [23] ), .B2(_01856_ ), .ZN(_03016_ ) );
NOR2_X1 _10270_ ( .A1(_03016_ ), .A2(_01833_ ), .ZN(_03017_ ) );
NAND3_X1 _10271_ ( .A1(_01578_ ), .A2(\u_csr.csr[1][23] ), .A3(_01579_ ), .ZN(_03018_ ) );
NAND4_X1 _10272_ ( .A1(_01584_ ), .A2(\u_csr.csr[2][23] ), .A3(_01590_ ), .A4(_01592_ ), .ZN(_03019_ ) );
NAND3_X1 _10273_ ( .A1(_01459_ ), .A2(\u_csr.csr[0][23] ), .A3(_01462_ ), .ZN(_03020_ ) );
AND2_X1 _10274_ ( .A1(_03019_ ), .A2(_03020_ ), .ZN(_03021_ ) );
AOI21_X1 _10275_ ( .A(_02492_ ), .B1(_03018_ ), .B2(_03021_ ), .ZN(_03022_ ) );
AOI211_X1 _10276_ ( .A(_01441_ ), .B(_02673_ ), .C1(_00847_ ), .C2(_00848_ ), .ZN(_03023_ ) );
NOR2_X1 _10277_ ( .A1(_03022_ ), .A2(_03023_ ), .ZN(_03024_ ) );
INV_X1 _10278_ ( .A(\de_pc [23] ), .ZN(_03025_ ) );
OAI22_X1 _10279_ ( .A1(_03024_ ), .A2(_01843_ ), .B1(_03025_ ), .B2(_01845_ ), .ZN(_03026_ ) );
OAI21_X1 _10280_ ( .A(_01070_ ), .B1(_03017_ ), .B2(_03026_ ), .ZN(_03027_ ) );
NOR2_X1 _10281_ ( .A1(_03016_ ), .A2(_01848_ ), .ZN(_03028_ ) );
NAND3_X1 _10282_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [23] ), .A3(_01512_ ), .ZN(_03029_ ) );
AND3_X1 _10283_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_03029_ ), .ZN(_03030_ ) );
OAI22_X1 _10284_ ( .A1(_01849_ ), .A2(_03025_ ), .B1(_01509_ ), .B2(_03030_ ), .ZN(_03031_ ) );
OAI21_X1 _10285_ ( .A(_00302_ ), .B1(_03028_ ), .B2(_03031_ ), .ZN(_03032_ ) );
NAND2_X1 _10286_ ( .A1(_03027_ ), .A2(_03032_ ), .ZN(_00159_ ) );
AND3_X1 _10287_ ( .A1(\ea_mask [0] ), .A2(\u_exu.eopt [15] ), .A3(\u_exu.ecsr [22] ), .ZN(_03033_ ) );
AOI211_X1 _10288_ ( .A(\u_arbiter.rvalid ), .B(_03033_ ), .C1(\ea_addr [22] ), .C2(_01521_ ), .ZN(_03034_ ) );
AOI21_X1 _10289_ ( .A(_01276_ ), .B1(_01998_ ), .B2(_02002_ ), .ZN(_03035_ ) );
NAND3_X1 _10290_ ( .A1(_01528_ ), .A2(_01143_ ), .A3(_01531_ ), .ZN(_03036_ ) );
AOI21_X1 _10291_ ( .A(_03035_ ), .B1(_01277_ ), .B2(_03036_ ), .ZN(_03037_ ) );
AOI21_X2 _10292_ ( .A(_01523_ ), .B1(\io_master_arsize [1] ), .B2(_03037_ ), .ZN(_03038_ ) );
AOI21_X2 _10293_ ( .A(_03034_ ), .B1(_03038_ ), .B2(\u_arbiter.rvalid ), .ZN(\ar_data [22] ) );
OR2_X2 _10294_ ( .A1(\ar_data [22] ), .A2(_01313_ ), .ZN(_03039_ ) );
AND3_X1 _10295_ ( .A1(_01307_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00938_ ), .ZN(_03040_ ) );
AOI221_X4 _10296_ ( .A(_03040_ ), .B1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00965_ ), .C1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(_01017_ ), .ZN(_03041_ ) );
NAND3_X1 _10297_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01547_ ), .ZN(_03042_ ) );
NAND3_X1 _10298_ ( .A1(_03041_ ), .A2(_01558_ ), .A3(_03042_ ), .ZN(_03043_ ) );
AOI22_X1 _10299_ ( .A1(_01322_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01752_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03044_ ) );
AOI21_X1 _10300_ ( .A(_01026_ ), .B1(_01542_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03045_ ) );
INV_X1 _10301_ ( .A(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03046_ ) );
OAI211_X1 _10302_ ( .A(_03044_ ), .B(_03045_ ), .C1(_03046_ ), .C2(_02403_ ), .ZN(_03047_ ) );
NAND3_X1 _10303_ ( .A1(_03043_ ), .A2(_01366_ ), .A3(_03047_ ), .ZN(_03048_ ) );
NAND3_X1 _10304_ ( .A1(_01292_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_01342_ ), .ZN(_03049_ ) );
NAND3_X1 _10305_ ( .A1(_01307_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01337_ ), .ZN(_03050_ ) );
NAND2_X1 _10306_ ( .A1(_03049_ ), .A2(_03050_ ), .ZN(_03051_ ) );
NAND3_X1 _10307_ ( .A1(_01292_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01337_ ), .ZN(_03052_ ) );
NAND2_X1 _10308_ ( .A1(_03052_ ), .A2(_01324_ ), .ZN(_03053_ ) );
AOI211_X1 _10309_ ( .A(_03051_ ), .B(_03053_ ), .C1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_01537_ ), .ZN(_03054_ ) );
OR2_X1 _10310_ ( .A1(_03054_ ), .A2(_01705_ ), .ZN(_03055_ ) );
NAND3_X1 _10311_ ( .A1(_01964_ ), .A2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(_01547_ ), .ZN(_03056_ ) );
AOI21_X1 _10312_ ( .A(_01345_ ), .B1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_01816_ ), .ZN(_03057_ ) );
INV_X1 _10313_ ( .A(\u_reg.rf[1][22] ), .ZN(_03058_ ) );
AOI21_X1 _10314_ ( .A(_03058_ ), .B1(_00936_ ), .B2(_00937_ ), .ZN(_03059_ ) );
OAI21_X1 _10315_ ( .A(_03056_ ), .B1(_03057_ ), .B2(_03059_ ), .ZN(_03060_ ) );
NOR2_X1 _10316_ ( .A1(_03060_ ), .A2(_01809_ ), .ZN(_03061_ ) );
OAI21_X1 _10317_ ( .A(_03048_ ), .B1(_03055_ ), .B2(_03061_ ), .ZN(_03062_ ) );
AOI21_X1 _10318_ ( .A(_01316_ ), .B1(_01536_ ), .B2(_03062_ ), .ZN(_03063_ ) );
NAND3_X1 _10319_ ( .A1(_03039_ ), .A2(_01370_ ), .A3(_03063_ ), .ZN(_03064_ ) );
NAND4_X1 _10320_ ( .A1(_01651_ ), .A2(\u_csr.csr[2][22] ), .A3(_01648_ ), .A4(_01649_ ), .ZN(_03065_ ) );
NAND3_X1 _10321_ ( .A1(_01577_ ), .A2(\u_csr.csr[1][22] ), .A3(_01651_ ), .ZN(_03066_ ) );
NAND4_X1 _10322_ ( .A1(_01653_ ), .A2(\u_csr.csr[0][22] ), .A3(_01654_ ), .A4(_01655_ ), .ZN(_03067_ ) );
NAND4_X1 _10323_ ( .A1(_01646_ ), .A2(_03065_ ), .A3(_03066_ ), .A4(_03067_ ), .ZN(_03068_ ) );
NAND2_X1 _10324_ ( .A1(_01575_ ), .A2(_03068_ ), .ZN(_03069_ ) );
NAND4_X1 _10325_ ( .A1(_01472_ ), .A2(_00850_ ), .A3(_00849_ ), .A4(_01443_ ), .ZN(_03070_ ) );
AOI21_X1 _10326_ ( .A(_01374_ ), .B1(_03069_ ), .B2(_03070_ ), .ZN(_03071_ ) );
AOI221_X4 _10327_ ( .A(_03071_ ), .B1(\de_pc [22] ), .B2(_01479_ ), .C1(_01105_ ), .C2(_01108_ ), .ZN(_03072_ ) );
NAND3_X1 _10328_ ( .A1(_03039_ ), .A2(_01484_ ), .A3(_03063_ ), .ZN(_03073_ ) );
NAND3_X1 _10329_ ( .A1(_01511_ ), .A2(\u_idu.imm_auipc_lui [22] ), .A3(_01512_ ), .ZN(_03074_ ) );
AND3_X1 _10330_ ( .A1(_01510_ ), .A2(_01517_ ), .A3(_03074_ ), .ZN(_03075_ ) );
NOR2_X1 _10331_ ( .A1(_01509_ ), .A2(_03075_ ), .ZN(_03076_ ) );
AOI211_X1 _10332_ ( .A(_03076_ ), .B(_01057_ ), .C1(\de_pc [22] ), .C2(_01492_ ), .ZN(_03077_ ) );
AOI221_X1 _10333_ ( .A(_02275_ ), .B1(_03064_ ), .B2(_03072_ ), .C1(_03073_ ), .C2(_03077_ ), .ZN(_00160_ ) );
NOR2_X1 _10334_ ( .A1(\u_exu.alu_ctrl [5] ), .A2(\u_exu.alu_ctrl [4] ), .ZN(_03078_ ) );
AND2_X1 _10335_ ( .A1(_03078_ ), .A2(fanout_net_19 ), .ZN(_03079_ ) );
INV_X1 _10336_ ( .A(_03079_ ), .ZN(_03080_ ) );
INV_X32 _10337_ ( .A(\u_exu.alu_ctrl [3] ), .ZN(_03081_ ) );
BUF_X32 _10338_ ( .A(_03081_ ), .Z(_03082_ ) );
BUF_X32 _10339_ ( .A(_03082_ ), .Z(_03083_ ) );
BUF_X16 _10340_ ( .A(_03083_ ), .Z(_03084_ ) );
AND3_X1 _10341_ ( .A1(_03084_ ), .A2(fanout_net_12 ), .A3(\u_exu.alu_p1 [0] ), .ZN(_03085_ ) );
INV_X1 _10342_ ( .A(\u_exu.alu_ctrl [4] ), .ZN(_03086_ ) );
NOR2_X1 _10343_ ( .A1(_03086_ ), .A2(\u_exu.alu_ctrl [5] ), .ZN(_03087_ ) );
INV_X1 _10344_ ( .A(fanout_net_12 ), .ZN(_03088_ ) );
CLKBUF_X2 _10345_ ( .A(_03088_ ), .Z(_03089_ ) );
NOR2_X1 _10346_ ( .A1(_03089_ ), .A2(\u_exu.alu_ctrl [3] ), .ZN(_03090_ ) );
OAI211_X1 _10347_ ( .A(fanout_net_19 ), .B(_03087_ ), .C1(_03090_ ), .C2(\u_exu.alu_p1 [0] ), .ZN(_03091_ ) );
AND2_X1 _10348_ ( .A1(\u_exu.alu_ctrl [5] ), .A2(\u_exu.alu_ctrl [4] ), .ZN(_03092_ ) );
AND2_X1 _10349_ ( .A1(_03092_ ), .A2(fanout_net_19 ), .ZN(_03093_ ) );
INV_X1 _10350_ ( .A(\u_exu.alu_p1 [0] ), .ZN(_03094_ ) );
NOR2_X1 _10351_ ( .A1(_03094_ ), .A2(fanout_net_12 ), .ZN(_03095_ ) );
INV_X1 _10352_ ( .A(fanout_net_14 ), .ZN(_03096_ ) );
AND2_X1 _10353_ ( .A1(_03095_ ), .A2(_03096_ ), .ZN(_03097_ ) );
INV_X1 _10354_ ( .A(\u_exu.alu_p2 [4] ), .ZN(_03098_ ) );
INV_X2 _10355_ ( .A(fanout_net_18 ), .ZN(_03099_ ) );
INV_X1 _10356_ ( .A(fanout_net_16 ), .ZN(_03100_ ) );
BUF_X4 _10357_ ( .A(_03100_ ), .Z(_03101_ ) );
BUF_X4 _10358_ ( .A(_03101_ ), .Z(_03102_ ) );
NAND4_X1 _10359_ ( .A1(_03097_ ), .A2(_03098_ ), .A3(_03099_ ), .A4(_03102_ ), .ZN(_03103_ ) );
AND2_X1 _10360_ ( .A1(_03078_ ), .A2(\u_exu.alu_ctrl [6] ), .ZN(_03104_ ) );
AOI21_X1 _10361_ ( .A(_03093_ ), .B1(_03103_ ), .B2(_03104_ ), .ZN(_03105_ ) );
XOR2_X1 _10362_ ( .A(fanout_net_12 ), .B(\u_exu.alu_p1 [0] ), .Z(_03106_ ) );
XOR2_X1 _10363_ ( .A(\u_exu.alu_p1 [6] ), .B(\u_exu.alu_p2 [6] ), .Z(_03107_ ) );
XOR2_X1 _10364_ ( .A(fanout_net_18 ), .B(\u_exu.alu_p1 [3] ), .Z(_03108_ ) );
XOR2_X1 _10365_ ( .A(\u_exu.alu_p1 [5] ), .B(\u_exu.alu_p2 [5] ), .Z(_03109_ ) );
NOR4_X1 _10366_ ( .A1(_03106_ ), .A2(_03107_ ), .A3(_03108_ ), .A4(_03109_ ), .ZN(_03110_ ) );
XOR2_X1 _10367_ ( .A(\u_exu.alu_p1 [23] ), .B(\u_exu.alu_p2 [23] ), .Z(_03111_ ) );
XOR2_X1 _10368_ ( .A(\u_exu.alu_p2 [17] ), .B(\u_exu.alu_p1 [17] ), .Z(_03112_ ) );
XOR2_X1 _10369_ ( .A(\u_exu.alu_p1 [18] ), .B(\u_exu.alu_p2 [18] ), .Z(_03113_ ) );
XOR2_X1 _10370_ ( .A(\u_exu.alu_p1 [21] ), .B(\u_exu.alu_p2 [21] ), .Z(_03114_ ) );
NOR4_X1 _10371_ ( .A1(_03111_ ), .A2(_03112_ ), .A3(_03113_ ), .A4(_03114_ ), .ZN(_03115_ ) );
XOR2_X1 _10372_ ( .A(\u_exu.alu_p1 [11] ), .B(\u_exu.alu_p2 [11] ), .Z(_03116_ ) );
XOR2_X1 _10373_ ( .A(\u_exu.alu_p1 [8] ), .B(\u_exu.alu_p2 [8] ), .Z(_03117_ ) );
XOR2_X1 _10374_ ( .A(\u_exu.alu_p1 [14] ), .B(\u_exu.alu_p2 [14] ), .Z(_03118_ ) );
XOR2_X1 _10375_ ( .A(\u_exu.alu_p1 [13] ), .B(\u_exu.alu_p2 [13] ), .Z(_03119_ ) );
NOR4_X1 _10376_ ( .A1(_03116_ ), .A2(_03117_ ), .A3(_03118_ ), .A4(_03119_ ), .ZN(_03120_ ) );
XOR2_X1 _10377_ ( .A(\u_exu.alu_p1 [30] ), .B(\u_exu.alu_p2 [30] ), .Z(_03121_ ) );
XOR2_X1 _10378_ ( .A(\u_exu.alu_p1 [27] ), .B(\u_exu.alu_p2 [27] ), .Z(_03122_ ) );
XOR2_X1 _10379_ ( .A(\u_exu.alu_p1 [29] ), .B(\u_exu.alu_p2 [29] ), .Z(_03123_ ) );
XOR2_X1 _10380_ ( .A(\u_exu.alu_p1 [24] ), .B(\u_exu.alu_p2 [24] ), .Z(_03124_ ) );
NOR4_X1 _10381_ ( .A1(_03121_ ), .A2(_03122_ ), .A3(_03123_ ), .A4(_03124_ ), .ZN(_03125_ ) );
AND4_X1 _10382_ ( .A1(_03110_ ), .A2(_03115_ ), .A3(_03120_ ), .A4(_03125_ ), .ZN(_03126_ ) );
XOR2_X1 _10383_ ( .A(\u_exu.alu_p2 [4] ), .B(\u_exu.alu_p1 [4] ), .Z(_03127_ ) );
XOR2_X1 _10384_ ( .A(fanout_net_14 ), .B(\u_exu.alu_p1 [1] ), .Z(_03128_ ) );
XOR2_X1 _10385_ ( .A(fanout_net_16 ), .B(\u_exu.alu_p1 [2] ), .Z(_03129_ ) );
AND2_X1 _10386_ ( .A1(\u_exu.alu_p1 [7] ), .A2(\u_exu.alu_p2 [7] ), .ZN(_03130_ ) );
NOR2_X1 _10387_ ( .A1(\u_exu.alu_p1 [7] ), .A2(\u_exu.alu_p2 [7] ), .ZN(_03131_ ) );
NOR2_X1 _10388_ ( .A1(_03130_ ), .A2(_03131_ ), .ZN(_03132_ ) );
NOR4_X1 _10389_ ( .A1(_03127_ ), .A2(_03128_ ), .A3(_03129_ ), .A4(_03132_ ), .ZN(_03133_ ) );
XOR2_X1 _10390_ ( .A(\u_exu.alu_p1 [12] ), .B(\u_exu.alu_p2 [12] ), .Z(_03134_ ) );
XOR2_X1 _10391_ ( .A(\u_exu.alu_p1 [10] ), .B(\u_exu.alu_p2 [10] ), .Z(_03135_ ) );
XOR2_X1 _10392_ ( .A(\u_exu.alu_p1 [15] ), .B(\u_exu.alu_p2 [15] ), .Z(_03136_ ) );
AND2_X1 _10393_ ( .A1(\u_exu.alu_p2 [9] ), .A2(\u_exu.alu_p1 [9] ), .ZN(_03137_ ) );
NOR2_X1 _10394_ ( .A1(\u_exu.alu_p2 [9] ), .A2(\u_exu.alu_p1 [9] ), .ZN(_03138_ ) );
NOR2_X1 _10395_ ( .A1(_03137_ ), .A2(_03138_ ), .ZN(_03139_ ) );
NOR4_X1 _10396_ ( .A1(_03134_ ), .A2(_03135_ ), .A3(_03136_ ), .A4(_03139_ ), .ZN(_03140_ ) );
XOR2_X1 _10397_ ( .A(\u_exu.alu_p1 [26] ), .B(\u_exu.alu_p2 [26] ), .Z(_03141_ ) );
XOR2_X1 _10398_ ( .A(\u_exu.alu_p1 [31] ), .B(\u_exu.alu_p2 [31] ), .Z(_03142_ ) );
AND2_X1 _10399_ ( .A1(\u_exu.alu_p1 [28] ), .A2(\u_exu.alu_p2 [28] ), .ZN(_03143_ ) );
NOR2_X1 _10400_ ( .A1(\u_exu.alu_p1 [28] ), .A2(\u_exu.alu_p2 [28] ), .ZN(_03144_ ) );
NOR2_X1 _10401_ ( .A1(_03143_ ), .A2(_03144_ ), .ZN(_03145_ ) );
AND2_X1 _10402_ ( .A1(\u_exu.alu_p1 [25] ), .A2(\u_exu.alu_p2 [25] ), .ZN(_03146_ ) );
NOR2_X1 _10403_ ( .A1(\u_exu.alu_p1 [25] ), .A2(\u_exu.alu_p2 [25] ), .ZN(_03147_ ) );
NOR2_X1 _10404_ ( .A1(_03146_ ), .A2(_03147_ ), .ZN(_03148_ ) );
NOR4_X1 _10405_ ( .A1(_03141_ ), .A2(_03142_ ), .A3(_03145_ ), .A4(_03148_ ), .ZN(_03149_ ) );
NOR2_X1 _10406_ ( .A1(\u_exu.alu_p1 [19] ), .A2(\u_exu.alu_p2 [19] ), .ZN(_03150_ ) );
AND2_X1 _10407_ ( .A1(\u_exu.alu_p1 [19] ), .A2(\u_exu.alu_p2 [19] ), .ZN(_03151_ ) );
AND2_X1 _10408_ ( .A1(\u_exu.alu_p1 [16] ), .A2(\u_exu.alu_p2 [16] ), .ZN(_03152_ ) );
NOR2_X1 _10409_ ( .A1(\u_exu.alu_p1 [16] ), .A2(\u_exu.alu_p2 [16] ), .ZN(_03153_ ) );
OAI22_X1 _10410_ ( .A1(_03150_ ), .A2(_03151_ ), .B1(_03152_ ), .B2(_03153_ ), .ZN(_03154_ ) );
XOR2_X1 _10411_ ( .A(\u_exu.alu_p1 [20] ), .B(\u_exu.alu_p2 [20] ), .Z(_03155_ ) );
AND2_X1 _10412_ ( .A1(\u_exu.alu_p1 [22] ), .A2(\u_exu.alu_p2 [22] ), .ZN(_03156_ ) );
NOR2_X1 _10413_ ( .A1(\u_exu.alu_p1 [22] ), .A2(\u_exu.alu_p2 [22] ), .ZN(_03157_ ) );
NOR2_X1 _10414_ ( .A1(_03156_ ), .A2(_03157_ ), .ZN(_03158_ ) );
NOR3_X1 _10415_ ( .A1(_03154_ ), .A2(_03155_ ), .A3(_03158_ ), .ZN(_03159_ ) );
AND4_X1 _10416_ ( .A1(_03133_ ), .A2(_03140_ ), .A3(_03149_ ), .A4(_03159_ ), .ZN(_03160_ ) );
NAND3_X1 _10417_ ( .A1(_03126_ ), .A2(_03160_ ), .A3(\u_exu.alu_ctrl [2] ), .ZN(_03161_ ) );
AND3_X1 _10418_ ( .A1(\u_exu.alu_ctrl [6] ), .A2(\u_exu.alu_ctrl [5] ), .A3(\u_exu.alu_ctrl [4] ), .ZN(_03162_ ) );
AND2_X1 _10419_ ( .A1(_03161_ ), .A2(_03162_ ), .ZN(_03163_ ) );
AND2_X1 _10420_ ( .A1(_03126_ ), .A2(_03160_ ), .ZN(_03164_ ) );
OAI21_X1 _10421_ ( .A(_03163_ ), .B1(\u_exu.alu_ctrl [2] ), .B2(_03164_ ), .ZN(_03165_ ) );
NAND2_X1 _10422_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [30] ), .ZN(_03166_ ) );
INV_X32 _10423_ ( .A(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03167_ ) );
BUF_X32 _10424_ ( .A(_03167_ ), .Z(_03168_ ) );
BUF_X32 _10425_ ( .A(_03168_ ), .Z(_03169_ ) );
BUF_X32 _10426_ ( .A(_03169_ ), .Z(_03170_ ) );
XNOR2_X1 _10427_ ( .A(_03166_ ), .B(_03170_ ), .ZN(_03171_ ) );
AND2_X1 _10428_ ( .A1(_03171_ ), .A2(\u_exu.alu_p1 [30] ), .ZN(_03172_ ) );
NAND2_X1 _10429_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [31] ), .ZN(_03173_ ) );
XNOR2_X1 _10430_ ( .A(_03173_ ), .B(_03170_ ), .ZN(_03174_ ) );
NAND2_X1 _10431_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [29] ), .ZN(_03175_ ) );
XNOR2_X1 _10432_ ( .A(_03175_ ), .B(_03170_ ), .ZN(_03176_ ) );
INV_X1 _10433_ ( .A(\u_exu.alu_p1 [29] ), .ZN(_03177_ ) );
XNOR2_X1 _10434_ ( .A(_03176_ ), .B(_03177_ ), .ZN(_03178_ ) );
INV_X1 _10435_ ( .A(_03178_ ), .ZN(_03179_ ) );
NAND2_X1 _10436_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [28] ), .ZN(_03180_ ) );
XNOR2_X1 _10437_ ( .A(_03180_ ), .B(_03170_ ), .ZN(_03181_ ) );
INV_X1 _10438_ ( .A(\u_exu.alu_p1 [28] ), .ZN(_03182_ ) );
XNOR2_X1 _10439_ ( .A(_03181_ ), .B(_03182_ ), .ZN(_03183_ ) );
INV_X1 _10440_ ( .A(_03183_ ), .ZN(_03184_ ) );
NAND2_X1 _10441_ ( .A1(_03081_ ), .A2(\u_exu.alu_p2 [15] ), .ZN(_03185_ ) );
XNOR2_X2 _10442_ ( .A(_03185_ ), .B(_03168_ ), .ZN(_03186_ ) );
XNOR2_X2 _10443_ ( .A(_03186_ ), .B(\u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03187_ ) );
NAND2_X4 _10444_ ( .A1(_03082_ ), .A2(\u_exu.alu_p2 [14] ), .ZN(_03188_ ) );
XNOR2_X2 _10445_ ( .A(_03188_ ), .B(_03168_ ), .ZN(_03189_ ) );
AND2_X1 _10446_ ( .A1(_03189_ ), .A2(\u_exu.alu_p1 [14] ), .ZN(_03190_ ) );
AND2_X1 _10447_ ( .A1(_03187_ ), .A2(_03190_ ), .ZN(_03191_ ) );
NAND2_X4 _10448_ ( .A1(_03081_ ), .A2(\u_exu.alu_p2 [9] ), .ZN(_03192_ ) );
XNOR2_X2 _10449_ ( .A(_03192_ ), .B(_03167_ ), .ZN(_03193_ ) );
XNOR2_X2 _10450_ ( .A(_03193_ ), .B(\u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03194_ ) );
NAND2_X1 _10451_ ( .A1(_03081_ ), .A2(\u_exu.alu_p2 [8] ), .ZN(_03195_ ) );
XNOR2_X2 _10452_ ( .A(_03195_ ), .B(_03168_ ), .ZN(_03196_ ) );
AND2_X4 _10453_ ( .A1(_03196_ ), .A2(\u_exu.alu_p1 [8] ), .ZN(_03197_ ) );
AND2_X4 _10454_ ( .A1(_03194_ ), .A2(_03197_ ), .ZN(_03198_ ) );
INV_X1 _10455_ ( .A(\u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03199_ ) );
AOI21_X2 _10456_ ( .A(_03198_ ), .B1(_03199_ ), .B2(_03193_ ), .ZN(_03200_ ) );
NAND2_X1 _10457_ ( .A1(_03081_ ), .A2(\u_exu.alu_p2 [10] ), .ZN(_03201_ ) );
XNOR2_X2 _10458_ ( .A(_03201_ ), .B(_03168_ ), .ZN(_03202_ ) );
INV_X1 _10459_ ( .A(\u_exu.alu_p1 [10] ), .ZN(_03203_ ) );
XNOR2_X1 _10460_ ( .A(_03202_ ), .B(_03203_ ), .ZN(_03204_ ) );
INV_X2 _10461_ ( .A(_03204_ ), .ZN(_03205_ ) );
NAND2_X4 _10462_ ( .A1(_03082_ ), .A2(\u_exu.alu_p2 [11] ), .ZN(_03206_ ) );
XNOR2_X2 _10463_ ( .A(_03206_ ), .B(_03168_ ), .ZN(_03207_ ) );
INV_X1 _10464_ ( .A(\u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03208_ ) );
AND2_X2 _10465_ ( .A1(_03207_ ), .A2(_03208_ ), .ZN(_03209_ ) );
NOR2_X1 _10466_ ( .A1(_03207_ ), .A2(_03208_ ), .ZN(_03210_ ) );
NOR4_X4 _10467_ ( .A1(_03200_ ), .A2(_03205_ ), .A3(_03209_ ), .A4(_03210_ ), .ZN(_03211_ ) );
XNOR2_X1 _10468_ ( .A(_03207_ ), .B(\u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03212_ ) );
AND2_X1 _10469_ ( .A1(_03202_ ), .A2(\u_exu.alu_p1 [10] ), .ZN(_03213_ ) );
AND2_X1 _10470_ ( .A1(_03212_ ), .A2(_03213_ ), .ZN(_03214_ ) );
NOR3_X4 _10471_ ( .A1(_03211_ ), .A2(_03209_ ), .A3(_03214_ ), .ZN(_03215_ ) );
NAND2_X4 _10472_ ( .A1(_03082_ ), .A2(\u_exu.alu_p2 [12] ), .ZN(_03216_ ) );
XNOR2_X2 _10473_ ( .A(_03216_ ), .B(_03168_ ), .ZN(_03217_ ) );
INV_X1 _10474_ ( .A(\u_exu.alu_p1 [12] ), .ZN(_03218_ ) );
XNOR2_X2 _10475_ ( .A(_03217_ ), .B(_03218_ ), .ZN(_03219_ ) );
NAND2_X4 _10476_ ( .A1(_03081_ ), .A2(\u_exu.alu_p2 [13] ), .ZN(_03220_ ) );
XNOR2_X2 _10477_ ( .A(_03220_ ), .B(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03221_ ) );
XNOR2_X1 _10478_ ( .A(_03221_ ), .B(\u_exu.alu_p1 [13] ), .ZN(_03222_ ) );
AND2_X4 _10479_ ( .A1(_03219_ ), .A2(_03222_ ), .ZN(_03223_ ) );
INV_X2 _10480_ ( .A(\u_exu.alu_p1 [14] ), .ZN(_03224_ ) );
XNOR2_X2 _10481_ ( .A(_03189_ ), .B(_03224_ ), .ZN(_03225_ ) );
AND2_X2 _10482_ ( .A1(_03225_ ), .A2(_03187_ ), .ZN(_03226_ ) );
AND2_X1 _10483_ ( .A1(_03223_ ), .A2(_03226_ ), .ZN(_03227_ ) );
INV_X1 _10484_ ( .A(_03227_ ), .ZN(_03228_ ) );
NOR2_X2 _10485_ ( .A1(_03215_ ), .A2(_03228_ ), .ZN(_03229_ ) );
INV_X1 _10486_ ( .A(_03226_ ), .ZN(_03230_ ) );
INV_X1 _10487_ ( .A(\u_exu.alu_p1 [13] ), .ZN(_03231_ ) );
NOR2_X1 _10488_ ( .A1(_03221_ ), .A2(_03231_ ), .ZN(_03232_ ) );
INV_X1 _10489_ ( .A(_03232_ ), .ZN(_03233_ ) );
AND2_X1 _10490_ ( .A1(_03217_ ), .A2(\u_exu.alu_p1 [12] ), .ZN(_03234_ ) );
NAND2_X1 _10491_ ( .A1(_03222_ ), .A2(_03234_ ), .ZN(_03235_ ) );
AOI21_X4 _10492_ ( .A(_03230_ ), .B1(_03233_ ), .B2(_03235_ ), .ZN(_03236_ ) );
OR2_X4 _10493_ ( .A1(_03229_ ), .A2(_03236_ ), .ZN(_03237_ ) );
INV_X1 _10494_ ( .A(\u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03238_ ) );
AOI211_X2 _10495_ ( .A(_03191_ ), .B(_03237_ ), .C1(_03238_ ), .C2(_03186_ ), .ZN(_03239_ ) );
INV_X1 _10496_ ( .A(\u_exu.alu_p1 [8] ), .ZN(_03240_ ) );
XNOR2_X1 _10497_ ( .A(_03196_ ), .B(_03240_ ), .ZN(_03241_ ) );
AND2_X1 _10498_ ( .A1(_03241_ ), .A2(_03194_ ), .ZN(_03242_ ) );
AND3_X1 _10499_ ( .A1(_03242_ ), .A2(_03212_ ), .A3(_03204_ ), .ZN(_03243_ ) );
NAND2_X1 _10500_ ( .A1(_03082_ ), .A2(\u_exu.alu_p2 [6] ), .ZN(_03244_ ) );
XNOR2_X2 _10501_ ( .A(_03244_ ), .B(_03169_ ), .ZN(_03245_ ) );
INV_X2 _10502_ ( .A(\u_exu.alu_p1 [6] ), .ZN(_03246_ ) );
XNOR2_X2 _10503_ ( .A(_03245_ ), .B(_03246_ ), .ZN(_03247_ ) );
NAND2_X4 _10504_ ( .A1(_03082_ ), .A2(\u_exu.alu_p2 [7] ), .ZN(_03248_ ) );
XNOR2_X2 _10505_ ( .A(_03248_ ), .B(_03168_ ), .ZN(_03249_ ) );
XNOR2_X2 _10506_ ( .A(_03249_ ), .B(\u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03250_ ) );
AND2_X4 _10507_ ( .A1(_03247_ ), .A2(_03250_ ), .ZN(_03251_ ) );
INV_X2 _10508_ ( .A(_03251_ ), .ZN(_03252_ ) );
NAND2_X1 _10509_ ( .A1(_03082_ ), .A2(\u_exu.alu_p2 [4] ), .ZN(_03253_ ) );
XNOR2_X2 _10510_ ( .A(_03253_ ), .B(_03169_ ), .ZN(_03254_ ) );
INV_X1 _10511_ ( .A(\u_exu.alu_p1 [4] ), .ZN(_03255_ ) );
XNOR2_X2 _10512_ ( .A(_03254_ ), .B(_03255_ ), .ZN(_03256_ ) );
NAND2_X1 _10513_ ( .A1(_03082_ ), .A2(\u_exu.alu_p2 [5] ), .ZN(_03257_ ) );
XNOR2_X2 _10514_ ( .A(_03257_ ), .B(_03169_ ), .ZN(_03258_ ) );
XNOR2_X2 _10515_ ( .A(_03258_ ), .B(\u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03259_ ) );
AND2_X2 _10516_ ( .A1(_03256_ ), .A2(_03259_ ), .ZN(_03260_ ) );
INV_X4 _10517_ ( .A(_03260_ ), .ZN(_03261_ ) );
NAND2_X4 _10518_ ( .A1(_03082_ ), .A2(fanout_net_18 ), .ZN(_03262_ ) );
XNOR2_X2 _10519_ ( .A(_03262_ ), .B(_03168_ ), .ZN(_03263_ ) );
XNOR2_X2 _10520_ ( .A(_03263_ ), .B(\u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03264_ ) );
NOR2_X4 _10521_ ( .A1(\u_exu.alu_ctrl [3] ), .A2(fanout_net_16 ), .ZN(_03265_ ) );
XNOR2_X1 _10522_ ( .A(_03265_ ), .B(fanout_net_11 ), .ZN(_03266_ ) );
INV_X1 _10523_ ( .A(\u_exu.alu_p1 [2] ), .ZN(_03267_ ) );
XNOR2_X1 _10524_ ( .A(_03266_ ), .B(_03267_ ), .ZN(_03268_ ) );
NAND2_X4 _10525_ ( .A1(_03082_ ), .A2(fanout_net_14 ), .ZN(_03269_ ) );
XNOR2_X2 _10526_ ( .A(_03269_ ), .B(_03168_ ), .ZN(_03270_ ) );
XNOR2_X2 _10527_ ( .A(_03270_ ), .B(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ), .ZN(_03271_ ) );
NAND3_X1 _10528_ ( .A1(_03083_ ), .A2(fanout_net_12 ), .A3(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ), .ZN(_03272_ ) );
OAI21_X2 _10529_ ( .A(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .B1(_03088_ ), .B2(\u_exu.alu_ctrl [3] ), .ZN(_03273_ ) );
AND3_X1 _10530_ ( .A1(_03271_ ), .A2(_03272_ ), .A3(_03273_ ), .ZN(_03274_ ) );
INV_X1 _10531_ ( .A(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ), .ZN(_03275_ ) );
AND2_X1 _10532_ ( .A1(_03270_ ), .A2(_03275_ ), .ZN(_03276_ ) );
OAI211_X2 _10533_ ( .A(_03264_ ), .B(_03268_ ), .C1(_03274_ ), .C2(_03276_ ), .ZN(_03277_ ) );
AND2_X1 _10534_ ( .A1(_03266_ ), .A2(\u_exu.alu_p1 [2] ), .ZN(_03278_ ) );
AND2_X2 _10535_ ( .A1(_03264_ ), .A2(_03278_ ), .ZN(_03279_ ) );
INV_X1 _10536_ ( .A(\u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03280_ ) );
AOI21_X2 _10537_ ( .A(_03279_ ), .B1(_03280_ ), .B2(_03263_ ), .ZN(_03281_ ) );
AOI211_X2 _10538_ ( .A(_03252_ ), .B(_03261_ ), .C1(_03277_ ), .C2(_03281_ ), .ZN(_03282_ ) );
NAND3_X1 _10539_ ( .A1(_03250_ ), .A2(\u_exu.alu_p1 [6] ), .A3(_03245_ ), .ZN(_03283_ ) );
INV_X1 _10540_ ( .A(_03249_ ), .ZN(_03284_ ) );
INV_X1 _10541_ ( .A(\u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03285_ ) );
AND2_X1 _10542_ ( .A1(_03258_ ), .A2(_03285_ ), .ZN(_03286_ ) );
AND2_X1 _10543_ ( .A1(_03254_ ), .A2(\u_exu.alu_p1 [4] ), .ZN(_03287_ ) );
AOI21_X1 _10544_ ( .A(_03286_ ), .B1(_03259_ ), .B2(_03287_ ), .ZN(_03288_ ) );
OAI221_X4 _10545_ ( .A(_03283_ ), .B1(\u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B2(_03284_ ), .C1(_03252_ ), .C2(_03288_ ), .ZN(_03289_ ) );
OAI211_X1 _10546_ ( .A(_03227_ ), .B(_03243_ ), .C1(_03282_ ), .C2(_03289_ ), .ZN(_03290_ ) );
AND2_X2 _10547_ ( .A1(_03239_ ), .A2(_03290_ ), .ZN(_03291_ ) );
INV_X4 _10548_ ( .A(_03291_ ), .ZN(_03292_ ) );
NAND2_X4 _10549_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [23] ), .ZN(_03293_ ) );
XNOR2_X2 _10550_ ( .A(_03293_ ), .B(_03169_ ), .ZN(_03294_ ) );
INV_X1 _10551_ ( .A(\u_exu.alu_p1 [23] ), .ZN(_03295_ ) );
XNOR2_X2 _10552_ ( .A(_03294_ ), .B(_03295_ ), .ZN(_03296_ ) );
NAND2_X4 _10553_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [22] ), .ZN(_03297_ ) );
XNOR2_X2 _10554_ ( .A(_03297_ ), .B(_03169_ ), .ZN(_03298_ ) );
INV_X1 _10555_ ( .A(\u_exu.alu_p1 [22] ), .ZN(_03299_ ) );
XNOR2_X2 _10556_ ( .A(_03298_ ), .B(_03299_ ), .ZN(_03300_ ) );
AND2_X1 _10557_ ( .A1(_03296_ ), .A2(_03300_ ), .ZN(_03301_ ) );
NAND2_X4 _10558_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [20] ), .ZN(_03302_ ) );
XNOR2_X2 _10559_ ( .A(_03302_ ), .B(_03169_ ), .ZN(_03303_ ) );
INV_X1 _10560_ ( .A(\u_exu.alu_p1 [20] ), .ZN(_03304_ ) );
XNOR2_X1 _10561_ ( .A(_03303_ ), .B(_03304_ ), .ZN(_03305_ ) );
NAND2_X4 _10562_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [21] ), .ZN(_03306_ ) );
XNOR2_X2 _10563_ ( .A(_03306_ ), .B(_03169_ ), .ZN(_03307_ ) );
XNOR2_X2 _10564_ ( .A(_03307_ ), .B(\u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03308_ ) );
AND2_X2 _10565_ ( .A1(_03305_ ), .A2(_03308_ ), .ZN(_03309_ ) );
AND2_X1 _10566_ ( .A1(_03301_ ), .A2(_03309_ ), .ZN(_03310_ ) );
NAND2_X4 _10567_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [16] ), .ZN(_03311_ ) );
XNOR2_X2 _10568_ ( .A(_03311_ ), .B(_03169_ ), .ZN(_03312_ ) );
INV_X1 _10569_ ( .A(\u_exu.alu_p1 [16] ), .ZN(_03313_ ) );
XNOR2_X1 _10570_ ( .A(_03312_ ), .B(_03313_ ), .ZN(_03314_ ) );
NAND2_X4 _10571_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [17] ), .ZN(_03315_ ) );
XNOR2_X2 _10572_ ( .A(_03315_ ), .B(_03169_ ), .ZN(_03316_ ) );
XNOR2_X2 _10573_ ( .A(_03316_ ), .B(\u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03317_ ) );
AND2_X1 _10574_ ( .A1(_03314_ ), .A2(_03317_ ), .ZN(_03318_ ) );
NAND2_X2 _10575_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [19] ), .ZN(_03319_ ) );
XNOR2_X2 _10576_ ( .A(_03319_ ), .B(_03170_ ), .ZN(_03320_ ) );
XNOR2_X1 _10577_ ( .A(_03320_ ), .B(\u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03321_ ) );
NAND2_X2 _10578_ ( .A1(_03083_ ), .A2(\u_exu.alu_p2 [18] ), .ZN(_03322_ ) );
XNOR2_X2 _10579_ ( .A(_03322_ ), .B(_03170_ ), .ZN(_03323_ ) );
INV_X1 _10580_ ( .A(\u_exu.alu_p1 [18] ), .ZN(_03324_ ) );
XNOR2_X1 _10581_ ( .A(_03323_ ), .B(_03324_ ), .ZN(_03325_ ) );
AND3_X1 _10582_ ( .A1(_03318_ ), .A2(_03321_ ), .A3(_03325_ ), .ZN(_03326_ ) );
NAND3_X4 _10583_ ( .A1(_03292_ ), .A2(_03310_ ), .A3(_03326_ ), .ZN(_03327_ ) );
AND2_X2 _10584_ ( .A1(_03312_ ), .A2(\u_exu.alu_p1 [16] ), .ZN(_03328_ ) );
AND2_X4 _10585_ ( .A1(_03317_ ), .A2(_03328_ ), .ZN(_03329_ ) );
INV_X1 _10586_ ( .A(\u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03330_ ) );
AOI21_X2 _10587_ ( .A(_03329_ ), .B1(_03330_ ), .B2(_03316_ ), .ZN(_03331_ ) );
INV_X1 _10588_ ( .A(_03325_ ), .ZN(_03332_ ) );
INV_X1 _10589_ ( .A(\u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03333_ ) );
AND2_X1 _10590_ ( .A1(_03320_ ), .A2(_03333_ ), .ZN(_03334_ ) );
NOR2_X1 _10591_ ( .A1(_03320_ ), .A2(_03333_ ), .ZN(_03335_ ) );
NOR4_X4 _10592_ ( .A1(_03331_ ), .A2(_03332_ ), .A3(_03334_ ), .A4(_03335_ ), .ZN(_03336_ ) );
AND2_X1 _10593_ ( .A1(_03323_ ), .A2(\u_exu.alu_p1 [18] ), .ZN(_03337_ ) );
AND2_X1 _10594_ ( .A1(_03321_ ), .A2(_03337_ ), .ZN(_03338_ ) );
NOR3_X4 _10595_ ( .A1(_03336_ ), .A2(_03334_ ), .A3(_03338_ ), .ZN(_03339_ ) );
INV_X1 _10596_ ( .A(_03310_ ), .ZN(_03340_ ) );
INV_X1 _10597_ ( .A(_03301_ ), .ZN(_03341_ ) );
AND2_X2 _10598_ ( .A1(_03303_ ), .A2(\u_exu.alu_p1 [20] ), .ZN(_03342_ ) );
AND2_X1 _10599_ ( .A1(_03308_ ), .A2(_03342_ ), .ZN(_03343_ ) );
INV_X1 _10600_ ( .A(\u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03344_ ) );
AOI21_X1 _10601_ ( .A(_03343_ ), .B1(_03344_ ), .B2(_03307_ ), .ZN(_03345_ ) );
OAI22_X1 _10602_ ( .A1(_03339_ ), .A2(_03340_ ), .B1(_03341_ ), .B2(_03345_ ), .ZN(_03346_ ) );
AND2_X1 _10603_ ( .A1(_03294_ ), .A2(\u_exu.alu_p1 [23] ), .ZN(_03347_ ) );
AND2_X1 _10604_ ( .A1(_03298_ ), .A2(\u_exu.alu_p1 [22] ), .ZN(_03348_ ) );
AND2_X1 _10605_ ( .A1(_03296_ ), .A2(_03348_ ), .ZN(_03349_ ) );
NOR3_X4 _10606_ ( .A1(_03346_ ), .A2(_03347_ ), .A3(_03349_ ), .ZN(_03350_ ) );
AND2_X4 _10607_ ( .A1(_03327_ ), .A2(_03350_ ), .ZN(_03351_ ) );
INV_X4 _10608_ ( .A(_03351_ ), .ZN(_03352_ ) );
NAND2_X1 _10609_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [27] ), .ZN(_03353_ ) );
XNOR2_X2 _10610_ ( .A(_03353_ ), .B(_03170_ ), .ZN(_03354_ ) );
INV_X1 _10611_ ( .A(\u_exu.alu_p1 [27] ), .ZN(_03355_ ) );
XNOR2_X1 _10612_ ( .A(_03354_ ), .B(_03355_ ), .ZN(_03356_ ) );
NAND2_X1 _10613_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [26] ), .ZN(_03357_ ) );
XNOR2_X1 _10614_ ( .A(_03357_ ), .B(_03170_ ), .ZN(_03358_ ) );
INV_X1 _10615_ ( .A(\u_exu.alu_p1 [26] ), .ZN(_03359_ ) );
XNOR2_X1 _10616_ ( .A(_03358_ ), .B(_03359_ ), .ZN(_03360_ ) );
AND2_X1 _10617_ ( .A1(_03356_ ), .A2(_03360_ ), .ZN(_03361_ ) );
NAND2_X1 _10618_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [24] ), .ZN(_03362_ ) );
XNOR2_X1 _10619_ ( .A(_03362_ ), .B(_03170_ ), .ZN(_03363_ ) );
INV_X1 _10620_ ( .A(\u_exu.alu_p1 [24] ), .ZN(_03364_ ) );
XNOR2_X1 _10621_ ( .A(_03363_ ), .B(_03364_ ), .ZN(_03365_ ) );
NAND2_X1 _10622_ ( .A1(_03084_ ), .A2(\u_exu.alu_p2 [25] ), .ZN(_03366_ ) );
XNOR2_X1 _10623_ ( .A(_03366_ ), .B(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03367_ ) );
XNOR2_X1 _10624_ ( .A(_03367_ ), .B(\u_exu.alu_p1 [25] ), .ZN(_03368_ ) );
NAND4_X4 _10625_ ( .A1(_03352_ ), .A2(_03361_ ), .A3(_03365_ ), .A4(_03368_ ), .ZN(_03369_ ) );
INV_X1 _10626_ ( .A(\u_exu.alu_p1 [25] ), .ZN(_03370_ ) );
NOR2_X1 _10627_ ( .A1(_03367_ ), .A2(_03370_ ), .ZN(_03371_ ) );
INV_X1 _10628_ ( .A(_03371_ ), .ZN(_03372_ ) );
AND2_X1 _10629_ ( .A1(_03363_ ), .A2(\u_exu.alu_p1 [24] ), .ZN(_03373_ ) );
INV_X1 _10630_ ( .A(_03373_ ), .ZN(_03374_ ) );
AND2_X1 _10631_ ( .A1(_03367_ ), .A2(_03370_ ), .ZN(_03375_ ) );
OAI21_X1 _10632_ ( .A(_03372_ ), .B1(_03374_ ), .B2(_03375_ ), .ZN(_03376_ ) );
AND3_X1 _10633_ ( .A1(_03376_ ), .A2(_03356_ ), .A3(_03360_ ), .ZN(_03377_ ) );
AND2_X1 _10634_ ( .A1(_03354_ ), .A2(\u_exu.alu_p1 [27] ), .ZN(_03378_ ) );
AND2_X1 _10635_ ( .A1(_03358_ ), .A2(\u_exu.alu_p1 [26] ), .ZN(_03379_ ) );
AND2_X1 _10636_ ( .A1(_03356_ ), .A2(_03379_ ), .ZN(_03380_ ) );
NOR3_X4 _10637_ ( .A1(_03377_ ), .A2(_03378_ ), .A3(_03380_ ), .ZN(_03381_ ) );
AOI211_X2 _10638_ ( .A(_03179_ ), .B(_03184_ ), .C1(_03369_ ), .C2(_03381_ ), .ZN(_03382_ ) );
AND2_X1 _10639_ ( .A1(_03181_ ), .A2(\u_exu.alu_p1 [28] ), .ZN(_03383_ ) );
AND2_X1 _10640_ ( .A1(_03178_ ), .A2(_03383_ ), .ZN(_03384_ ) );
AOI21_X1 _10641_ ( .A(_03384_ ), .B1(\u_exu.alu_p1 [29] ), .B2(_03176_ ), .ZN(_03385_ ) );
INV_X1 _10642_ ( .A(_03385_ ), .ZN(_03386_ ) );
NOR2_X2 _10643_ ( .A1(_03382_ ), .A2(_03386_ ), .ZN(_03387_ ) );
INV_X2 _10644_ ( .A(_03387_ ), .ZN(_03388_ ) );
INV_X1 _10645_ ( .A(\u_exu.alu_p1 [30] ), .ZN(_03389_ ) );
XNOR2_X1 _10646_ ( .A(_03171_ ), .B(_03389_ ), .ZN(_03390_ ) );
AOI221_X1 _10647_ ( .A(_03172_ ), .B1(\u_exu.alu_p1 [31] ), .B2(_03174_ ), .C1(_03388_ ), .C2(_03390_ ), .ZN(_03391_ ) );
NOR2_X1 _10648_ ( .A1(_03174_ ), .A2(\u_exu.alu_p1 [31] ), .ZN(_03392_ ) );
OR3_X1 _10649_ ( .A1(_03391_ ), .A2(\u_exu.alu_ctrl [1] ), .A3(_03392_ ), .ZN(_03393_ ) );
AOI21_X2 _10650_ ( .A(_03172_ ), .B1(_03388_ ), .B2(_03390_ ), .ZN(_03394_ ) );
INV_X1 _10651_ ( .A(\u_exu.alu_p1 [31] ), .ZN(_03395_ ) );
XNOR2_X1 _10652_ ( .A(_03174_ ), .B(_03395_ ), .ZN(_03396_ ) );
NAND2_X1 _10653_ ( .A1(_03394_ ), .A2(_03396_ ), .ZN(_03397_ ) );
OAI211_X2 _10654_ ( .A(_03397_ ), .B(\u_exu.alu_ctrl [1] ), .C1(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ), .C2(_03396_ ), .ZN(_03398_ ) );
NAND3_X1 _10655_ ( .A1(_03393_ ), .A2(\u_exu.alu_ctrl [2] ), .A3(_03398_ ), .ZN(_03399_ ) );
INV_X1 _10656_ ( .A(\u_exu.alu_ctrl [5] ), .ZN(_03400_ ) );
NOR2_X2 _10657_ ( .A1(_03400_ ), .A2(\u_exu.alu_ctrl [4] ), .ZN(_03401_ ) );
NAND3_X1 _10658_ ( .A1(_03399_ ), .A2(\u_exu.alu_ctrl [6] ), .A3(_03401_ ), .ZN(_03402_ ) );
AOI21_X1 _10659_ ( .A(\u_exu.alu_ctrl [2] ), .B1(_03393_ ), .B2(_03398_ ), .ZN(_03403_ ) );
OAI21_X1 _10660_ ( .A(_03165_ ), .B1(_03402_ ), .B2(_03403_ ), .ZN(_03404_ ) );
NOR2_X1 _10661_ ( .A1(_03267_ ), .A2(fanout_net_12 ), .ZN(_03405_ ) );
AND2_X1 _10662_ ( .A1(fanout_net_12 ), .A2(\u_exu.alu_p1 [3] ), .ZN(_03406_ ) );
NOR2_X1 _10663_ ( .A1(_03405_ ), .A2(_03406_ ), .ZN(_03407_ ) );
NOR2_X1 _10664_ ( .A1(_03407_ ), .A2(_03096_ ), .ZN(_03408_ ) );
AND3_X1 _10665_ ( .A1(_03096_ ), .A2(fanout_net_12 ), .A3(\u_exu.alu_p1 [1] ), .ZN(_03409_ ) );
NOR4_X1 _10666_ ( .A1(_03408_ ), .A2(fanout_net_16 ), .A3(_03097_ ), .A4(_03409_ ), .ZN(_03410_ ) );
NOR2_X1 _10667_ ( .A1(_03255_ ), .A2(fanout_net_12 ), .ZN(_03411_ ) );
AND2_X1 _10668_ ( .A1(fanout_net_12 ), .A2(\u_exu.alu_p1 [5] ), .ZN(_03412_ ) );
OAI21_X1 _10669_ ( .A(_03096_ ), .B1(_03411_ ), .B2(_03412_ ), .ZN(_03413_ ) );
NOR2_X1 _10670_ ( .A1(_03246_ ), .A2(fanout_net_12 ), .ZN(_03414_ ) );
AND2_X1 _10671_ ( .A1(fanout_net_12 ), .A2(\u_exu.alu_p1 [7] ), .ZN(_03415_ ) );
OAI21_X1 _10672_ ( .A(fanout_net_14 ), .B1(_03414_ ), .B2(_03415_ ), .ZN(_03416_ ) );
AND2_X1 _10673_ ( .A1(_03413_ ), .A2(_03416_ ), .ZN(_03417_ ) );
AOI211_X1 _10674_ ( .A(fanout_net_18 ), .B(_03410_ ), .C1(fanout_net_16 ), .C2(_03417_ ), .ZN(_03418_ ) );
NOR2_X1 _10675_ ( .A1(_03203_ ), .A2(fanout_net_12 ), .ZN(_03419_ ) );
AND2_X1 _10676_ ( .A1(fanout_net_12 ), .A2(\u_exu.alu_p1 [11] ), .ZN(_03420_ ) );
OR3_X1 _10677_ ( .A1(_03419_ ), .A2(_03420_ ), .A3(_03096_ ), .ZN(_03421_ ) );
NOR2_X1 _10678_ ( .A1(_03240_ ), .A2(fanout_net_12 ), .ZN(_03422_ ) );
AND2_X1 _10679_ ( .A1(fanout_net_12 ), .A2(\u_exu.alu_p1 [9] ), .ZN(_03423_ ) );
OR3_X1 _10680_ ( .A1(_03422_ ), .A2(_03423_ ), .A3(fanout_net_14 ), .ZN(_03424_ ) );
NAND3_X1 _10681_ ( .A1(_03421_ ), .A2(_03424_ ), .A3(_03100_ ), .ZN(_03425_ ) );
NOR2_X1 _10682_ ( .A1(_03224_ ), .A2(fanout_net_12 ), .ZN(_03426_ ) );
AND2_X1 _10683_ ( .A1(\u_exu.alu_p1 [15] ), .A2(fanout_net_12 ), .ZN(_03427_ ) );
OR3_X1 _10684_ ( .A1(_03426_ ), .A2(_03427_ ), .A3(_03096_ ), .ZN(_03428_ ) );
NOR2_X1 _10685_ ( .A1(_03218_ ), .A2(fanout_net_12 ), .ZN(_03429_ ) );
AND2_X1 _10686_ ( .A1(\u_exu.alu_p1 [13] ), .A2(fanout_net_12 ), .ZN(_03430_ ) );
OR3_X1 _10687_ ( .A1(_03429_ ), .A2(_03430_ ), .A3(fanout_net_14 ), .ZN(_03431_ ) );
NAND3_X1 _10688_ ( .A1(_03428_ ), .A2(_03431_ ), .A3(fanout_net_16 ), .ZN(_03432_ ) );
AOI21_X1 _10689_ ( .A(_03099_ ), .B1(_03425_ ), .B2(_03432_ ), .ZN(_03433_ ) );
OR3_X1 _10690_ ( .A1(_03418_ ), .A2(\u_exu.alu_p2 [4] ), .A3(_03433_ ), .ZN(_03434_ ) );
INV_X1 _10691_ ( .A(fanout_net_19 ), .ZN(_03435_ ) );
AND2_X1 _10692_ ( .A1(_03087_ ), .A2(_03435_ ), .ZN(_03436_ ) );
INV_X2 _10693_ ( .A(_03436_ ), .ZN(_03437_ ) );
AOI21_X1 _10694_ ( .A(_03437_ ), .B1(\u_exu.alu_ctrl [1] ), .B2(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_Y_$_MUX__B_A_$_NOR__Y_A_$_ANDNOT__Y_B ), .ZN(_03438_ ) );
NAND2_X1 _10695_ ( .A1(_03434_ ), .A2(_03438_ ), .ZN(_03439_ ) );
NOR2_X1 _10696_ ( .A1(_03324_ ), .A2(fanout_net_12 ), .ZN(_03440_ ) );
AND2_X1 _10697_ ( .A1(\u_exu.alu_p1 [19] ), .A2(fanout_net_12 ), .ZN(_03441_ ) );
OR3_X1 _10698_ ( .A1(_03440_ ), .A2(_03441_ ), .A3(_03096_ ), .ZN(_03442_ ) );
NOR2_X1 _10699_ ( .A1(_03313_ ), .A2(fanout_net_12 ), .ZN(_03443_ ) );
AND2_X1 _10700_ ( .A1(\u_exu.alu_p1 [17] ), .A2(fanout_net_12 ), .ZN(_03444_ ) );
OR3_X1 _10701_ ( .A1(_03443_ ), .A2(_03444_ ), .A3(fanout_net_14 ), .ZN(_03445_ ) );
NAND2_X1 _10702_ ( .A1(_03442_ ), .A2(_03445_ ), .ZN(_03446_ ) );
NAND2_X1 _10703_ ( .A1(_03446_ ), .A2(_03100_ ), .ZN(_03447_ ) );
NOR2_X1 _10704_ ( .A1(_03304_ ), .A2(fanout_net_12 ), .ZN(_03448_ ) );
AND2_X1 _10705_ ( .A1(\u_exu.alu_p1 [21] ), .A2(fanout_net_12 ), .ZN(_03449_ ) );
OR3_X1 _10706_ ( .A1(_03448_ ), .A2(_03449_ ), .A3(fanout_net_14 ), .ZN(_03450_ ) );
AND2_X1 _10707_ ( .A1(fanout_net_12 ), .A2(\u_exu.alu_p1 [23] ), .ZN(_03451_ ) );
INV_X1 _10708_ ( .A(_03451_ ), .ZN(_03452_ ) );
OAI211_X1 _10709_ ( .A(_03452_ ), .B(fanout_net_14 ), .C1(fanout_net_12 ), .C2(_03299_ ), .ZN(_03453_ ) );
NAND2_X1 _10710_ ( .A1(_03450_ ), .A2(_03453_ ), .ZN(_03454_ ) );
NAND2_X1 _10711_ ( .A1(_03454_ ), .A2(fanout_net_16 ), .ZN(_03455_ ) );
AND3_X1 _10712_ ( .A1(_03447_ ), .A2(_03455_ ), .A3(_03099_ ), .ZN(_03456_ ) );
NOR2_X1 _10713_ ( .A1(_03182_ ), .A2(fanout_net_12 ), .ZN(_03457_ ) );
AND2_X1 _10714_ ( .A1(\u_exu.alu_p1 [29] ), .A2(fanout_net_12 ), .ZN(_03458_ ) );
NOR2_X1 _10715_ ( .A1(_03457_ ), .A2(_03458_ ), .ZN(_03459_ ) );
MUX2_X1 _10716_ ( .A(_03389_ ), .B(_03395_ ), .S(fanout_net_13 ), .Z(_03460_ ) );
MUX2_X1 _10717_ ( .A(_03459_ ), .B(_03460_ ), .S(fanout_net_14 ), .Z(_03461_ ) );
OR2_X1 _10718_ ( .A1(_03461_ ), .A2(_03100_ ), .ZN(_03462_ ) );
NOR2_X1 _10719_ ( .A1(_03359_ ), .A2(fanout_net_13 ), .ZN(_03463_ ) );
INV_X1 _10720_ ( .A(_03463_ ), .ZN(_03464_ ) );
AND2_X1 _10721_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [27] ), .ZN(_03465_ ) );
INV_X1 _10722_ ( .A(_03465_ ), .ZN(_03466_ ) );
NAND3_X1 _10723_ ( .A1(_03464_ ), .A2(fanout_net_14 ), .A3(_03466_ ), .ZN(_03467_ ) );
NOR2_X1 _10724_ ( .A1(_03364_ ), .A2(fanout_net_13 ), .ZN(_03468_ ) );
INV_X1 _10725_ ( .A(_03468_ ), .ZN(_03469_ ) );
BUF_X4 _10726_ ( .A(_03096_ ), .Z(_03470_ ) );
AND2_X1 _10727_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [25] ), .ZN(_03471_ ) );
INV_X1 _10728_ ( .A(_03471_ ), .ZN(_03472_ ) );
NAND3_X1 _10729_ ( .A1(_03469_ ), .A2(_03470_ ), .A3(_03472_ ), .ZN(_03473_ ) );
NAND2_X1 _10730_ ( .A1(_03467_ ), .A2(_03473_ ), .ZN(_03474_ ) );
OAI21_X1 _10731_ ( .A(_03462_ ), .B1(fanout_net_16 ), .B2(_03474_ ), .ZN(_03475_ ) );
AOI21_X1 _10732_ ( .A(_03456_ ), .B1(_03475_ ), .B2(fanout_net_18 ), .ZN(_03476_ ) );
AOI21_X1 _10733_ ( .A(_03439_ ), .B1(\u_exu.alu_p2 [4] ), .B2(_03476_ ), .ZN(_03477_ ) );
OR2_X1 _10734_ ( .A1(_03477_ ), .A2(_03104_ ), .ZN(_03478_ ) );
OAI21_X1 _10735_ ( .A(_03105_ ), .B1(_03404_ ), .B2(_03478_ ), .ZN(_03479_ ) );
AND2_X1 _10736_ ( .A1(_03401_ ), .A2(fanout_net_19 ), .ZN(_03480_ ) );
INV_X1 _10737_ ( .A(_03480_ ), .ZN(_03481_ ) );
BUF_X4 _10738_ ( .A(_03093_ ), .Z(_03482_ ) );
NAND2_X1 _10739_ ( .A1(_03106_ ), .A2(_03482_ ), .ZN(_03483_ ) );
AND3_X2 _10740_ ( .A1(_03479_ ), .A2(_03481_ ), .A3(_03483_ ), .ZN(_03484_ ) );
AND2_X1 _10741_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [0] ), .ZN(_03485_ ) );
INV_X1 _10742_ ( .A(_03485_ ), .ZN(_03486_ ) );
OAI21_X1 _10743_ ( .A(fanout_net_11 ), .B1(fanout_net_13 ), .B2(\u_exu.alu_p1 [0] ), .ZN(_03487_ ) );
AND3_X1 _10744_ ( .A1(_03480_ ), .A2(_03486_ ), .A3(_03487_ ), .ZN(_03488_ ) );
OAI221_X2 _10745_ ( .A(_03080_ ), .B1(_03085_ ), .B2(_03091_ ), .C1(_03484_ ), .C2(_03488_ ), .ZN(_03489_ ) );
BUF_X2 _10746_ ( .A(_03086_ ), .Z(_03490_ ) );
NAND4_X1 _10747_ ( .A1(_03400_ ), .A2(_03490_ ), .A3(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ), .A4(fanout_net_19 ), .ZN(_03491_ ) );
AND3_X4 _10748_ ( .A1(_03489_ ), .A2(_01475_ ), .A3(_03491_ ), .ZN(_03492_ ) );
BUF_X4 _10749_ ( .A(_00744_ ), .Z(_03493_ ) );
OR2_X4 _10750_ ( .A1(_03492_ ), .A2(_03493_ ), .ZN(_03494_ ) );
INV_X1 _10751_ ( .A(_01505_ ), .ZN(_03495_ ) );
AOI211_X1 _10752_ ( .A(_00892_ ), .B(_03495_ ), .C1(_01106_ ), .C2(_01109_ ), .ZN(_03496_ ) );
NAND2_X4 _10753_ ( .A1(_03494_ ), .A2(_03496_ ), .ZN(_03497_ ) );
BUF_X8 _10754_ ( .A(_03497_ ), .Z(_03498_ ) );
INV_X1 _10755_ ( .A(_01440_ ), .ZN(_03499_ ) );
BUF_X4 _10756_ ( .A(_03499_ ), .Z(_03500_ ) );
XNOR2_X1 _10757_ ( .A(_00928_ ), .B(_01295_ ), .ZN(_03501_ ) );
XNOR2_X1 _10758_ ( .A(_00989_ ), .B(_01304_ ), .ZN(_03502_ ) );
XNOR2_X1 _10759_ ( .A(_01049_ ), .B(_01289_ ), .ZN(_03503_ ) );
OR3_X1 _10760_ ( .A1(_00925_ ), .A2(_00888_ ), .A3(_01299_ ), .ZN(_03504_ ) );
NAND4_X1 _10761_ ( .A1(_03501_ ), .A2(_03502_ ), .A3(_03503_ ), .A4(_03504_ ), .ZN(_03505_ ) );
AOI21_X1 _10762_ ( .A(_03505_ ), .B1(_01028_ ), .B2(_01308_ ), .ZN(_03506_ ) );
AND2_X4 _10763_ ( .A1(_01286_ ), .A2(_03506_ ), .ZN(_03507_ ) );
INV_X4 _10764_ ( .A(_03507_ ), .ZN(_03508_ ) );
BUF_X16 _10765_ ( .A(_03508_ ), .Z(_03509_ ) );
BUF_X16 _10766_ ( .A(_03509_ ), .Z(_03510_ ) );
BUF_X16 _10767_ ( .A(_03510_ ), .Z(_03511_ ) );
NOR2_X1 _10768_ ( .A1(\ar_data [31] ), .A2(_03511_ ), .ZN(_03512_ ) );
NAND2_X1 _10769_ ( .A1(_00669_ ), .A2(_01078_ ), .ZN(_03513_ ) );
AOI21_X1 _10770_ ( .A(_00687_ ), .B1(_00692_ ), .B2(_00701_ ), .ZN(_03514_ ) );
AND2_X2 _10771_ ( .A1(_03513_ ), .A2(_03514_ ), .ZN(_03515_ ) );
INV_X1 _10772_ ( .A(_03515_ ), .ZN(_03516_ ) );
BUF_X4 _10773_ ( .A(_00955_ ), .Z(_03517_ ) );
BUF_X4 _10774_ ( .A(_03517_ ), .Z(_03518_ ) );
BUF_X2 _10775_ ( .A(_03518_ ), .Z(_03519_ ) );
BUF_X4 _10776_ ( .A(_00928_ ), .Z(_03520_ ) );
BUF_X4 _10777_ ( .A(_03520_ ), .Z(_03521_ ) );
BUF_X4 _10778_ ( .A(_03521_ ), .Z(_03522_ ) );
BUF_X2 _10779_ ( .A(_00749_ ), .Z(_03523_ ) );
BUF_X2 _10780_ ( .A(_03523_ ), .Z(_03524_ ) );
NAND3_X1 _10781_ ( .A1(_03522_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03525_ ) );
NAND3_X1 _10782_ ( .A1(_03522_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03526_ ) );
BUF_X2 _10783_ ( .A(_00989_ ), .Z(_03527_ ) );
BUF_X4 _10784_ ( .A(_03527_ ), .Z(_03528_ ) );
BUF_X4 _10785_ ( .A(_03528_ ), .Z(_03529_ ) );
NAND3_X1 _10786_ ( .A1(_03529_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03530_ ) );
NAND3_X1 _10787_ ( .A1(_03525_ ), .A2(_03526_ ), .A3(_03530_ ), .ZN(_03531_ ) );
BUF_X4 _10788_ ( .A(_01019_ ), .Z(_03532_ ) );
BUF_X4 _10789_ ( .A(_03532_ ), .Z(_03533_ ) );
BUF_X4 _10790_ ( .A(_03533_ ), .Z(_03534_ ) );
BUF_X4 _10791_ ( .A(_03534_ ), .Z(_03535_ ) );
AOI211_X1 _10792_ ( .A(_03519_ ), .B(_03531_ ), .C1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03535_ ), .ZN(_03536_ ) );
BUF_X4 _10793_ ( .A(_01028_ ), .Z(_03537_ ) );
CLKBUF_X2 _10794_ ( .A(_03537_ ), .Z(_03538_ ) );
BUF_X4 _10795_ ( .A(_01049_ ), .Z(_03539_ ) );
AOI21_X1 _10796_ ( .A(_03539_ ), .B1(_03534_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03540_ ) );
CLKBUF_X2 _10797_ ( .A(_03528_ ), .Z(_03541_ ) );
NAND3_X1 _10798_ ( .A1(_03541_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03542_ ) );
BUF_X2 _10799_ ( .A(_03523_ ), .Z(_03543_ ) );
NAND3_X1 _10800_ ( .A1(_03522_ ), .A2(_03543_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03544_ ) );
NAND3_X1 _10801_ ( .A1(_03541_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03545_ ) );
AND4_X1 _10802_ ( .A1(_03540_ ), .A2(_03542_ ), .A3(_03544_ ), .A4(_03545_ ), .ZN(_03546_ ) );
NOR3_X1 _10803_ ( .A1(_03536_ ), .A2(_03538_ ), .A3(_03546_ ), .ZN(_03547_ ) );
CLKBUF_X2 _10804_ ( .A(_00989_ ), .Z(_03548_ ) );
CLKBUF_X2 _10805_ ( .A(_03548_ ), .Z(_03549_ ) );
AND3_X1 _10806_ ( .A1(_03549_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03550_ ) );
BUF_X4 _10807_ ( .A(_03533_ ), .Z(_03551_ ) );
BUF_X4 _10808_ ( .A(_00980_ ), .Z(_03552_ ) );
BUF_X4 _10809_ ( .A(_03552_ ), .Z(_03553_ ) );
AOI221_X4 _10810_ ( .A(_03550_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03553_ ), .ZN(_03554_ ) );
BUF_X4 _10811_ ( .A(_01049_ ), .Z(_03555_ ) );
BUF_X4 _10812_ ( .A(_03555_ ), .Z(_03556_ ) );
BUF_X2 _10813_ ( .A(_03556_ ), .Z(_03557_ ) );
BUF_X4 _10814_ ( .A(_03522_ ), .Z(_03558_ ) );
BUF_X4 _10815_ ( .A(_03558_ ), .Z(_03559_ ) );
BUF_X2 _10816_ ( .A(_00749_ ), .Z(_03560_ ) );
BUF_X2 _10817_ ( .A(_03560_ ), .Z(_03561_ ) );
BUF_X4 _10818_ ( .A(_03561_ ), .Z(_03562_ ) );
BUF_X4 _10819_ ( .A(_03562_ ), .Z(_03563_ ) );
NAND3_X1 _10820_ ( .A1(_03559_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03564_ ) );
NAND3_X1 _10821_ ( .A1(_03554_ ), .A2(_03557_ ), .A3(_03564_ ), .ZN(_03565_ ) );
OR3_X1 _10822_ ( .A1(_00925_ ), .A2(_03561_ ), .A3(_01346_ ), .ZN(_03566_ ) );
BUF_X4 _10823_ ( .A(_00956_ ), .Z(_03567_ ) );
AOI21_X1 _10824_ ( .A(_03556_ ), .B1(_03566_ ), .B2(_03567_ ), .ZN(_03568_ ) );
BUF_X4 _10825_ ( .A(_03543_ ), .Z(_03569_ ) );
NAND3_X1 _10826_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03570_ ) );
BUF_X2 _10827_ ( .A(_03529_ ), .Z(_03571_ ) );
NAND3_X1 _10828_ ( .A1(_03571_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03572_ ) );
NAND3_X1 _10829_ ( .A1(_03568_ ), .A2(_03570_ ), .A3(_03572_ ), .ZN(_03573_ ) );
AND2_X1 _10830_ ( .A1(_03573_ ), .A2(_03538_ ), .ZN(_03574_ ) );
AOI21_X1 _10831_ ( .A(_03547_ ), .B1(_03565_ ), .B2(_03574_ ), .ZN(_03575_ ) );
OAI21_X1 _10832_ ( .A(_03516_ ), .B1(_03507_ ), .B2(_03575_ ), .ZN(_03576_ ) );
OAI21_X1 _10833_ ( .A(_03500_ ), .B1(_03512_ ), .B2(_03576_ ), .ZN(_03577_ ) );
NOR2_X1 _10834_ ( .A1(_01482_ ), .A2(_01490_ ), .ZN(_03578_ ) );
CLKBUF_X2 _10835_ ( .A(_01440_ ), .Z(_03579_ ) );
CLKBUF_X2 _10836_ ( .A(_03579_ ), .Z(_03580_ ) );
NAND3_X1 _10837_ ( .A1(_01470_ ), .A2(_03580_ ), .A3(_01473_ ), .ZN(_03581_ ) );
AND3_X1 _10838_ ( .A1(_03577_ ), .A2(_03578_ ), .A3(_03581_ ), .ZN(_03582_ ) );
AOI211_X1 _10839_ ( .A(_00860_ ), .B(_01493_ ), .C1(_00900_ ), .C2(_02359_ ), .ZN(_03583_ ) );
OAI21_X1 _10840_ ( .A(_00302_ ), .B1(_03582_ ), .B2(_03583_ ), .ZN(_03584_ ) );
NAND2_X1 _10841_ ( .A1(_03498_ ), .A2(_03584_ ), .ZN(_00161_ ) );
INV_X1 _10842_ ( .A(_03578_ ), .ZN(_03585_ ) );
BUF_X4 _10843_ ( .A(_03585_ ), .Z(_03586_ ) );
AND3_X1 _10844_ ( .A1(_01595_ ), .A2(_03580_ ), .A3(_01598_ ), .ZN(_03587_ ) );
NOR2_X2 _10845_ ( .A1(\ar_data [30] ), .A2(_03511_ ), .ZN(_03588_ ) );
AND3_X1 _10846_ ( .A1(_03528_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03589_ ) );
BUF_X4 _10847_ ( .A(_03520_ ), .Z(_03590_ ) );
AND3_X1 _10848_ ( .A1(_03590_ ), .A2(_03523_ ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03591_ ) );
AND3_X1 _10849_ ( .A1(_03548_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03592_ ) );
OR3_X1 _10850_ ( .A1(_03589_ ), .A2(_03591_ ), .A3(_03592_ ), .ZN(_03593_ ) );
AOI211_X1 _10851_ ( .A(_03519_ ), .B(_03593_ ), .C1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03535_ ), .ZN(_03594_ ) );
AOI21_X1 _10852_ ( .A(_03555_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03595_ ) );
NAND3_X1 _10853_ ( .A1(_03541_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03596_ ) );
NAND3_X1 _10854_ ( .A1(_03522_ ), .A2(_03543_ ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03597_ ) );
NAND3_X1 _10855_ ( .A1(_03541_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03598_ ) );
AND4_X1 _10856_ ( .A1(_03595_ ), .A2(_03596_ ), .A3(_03597_ ), .A4(_03598_ ), .ZN(_03599_ ) );
NOR3_X1 _10857_ ( .A1(_03594_ ), .A2(_03538_ ), .A3(_03599_ ), .ZN(_03600_ ) );
BUF_X4 _10858_ ( .A(_03556_ ), .Z(_03601_ ) );
OR3_X1 _10859_ ( .A1(_00925_ ), .A2(_03543_ ), .A3(_01552_ ), .ZN(_03602_ ) );
AOI21_X1 _10860_ ( .A(_03601_ ), .B1(_03602_ ), .B2(_03567_ ), .ZN(_03603_ ) );
NAND3_X1 _10861_ ( .A1(_03559_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03604_ ) );
BUF_X4 _10862_ ( .A(_03528_ ), .Z(_03605_ ) );
BUF_X4 _10863_ ( .A(_03605_ ), .Z(_03606_ ) );
BUF_X4 _10864_ ( .A(_03606_ ), .Z(_03607_ ) );
NAND3_X1 _10865_ ( .A1(_03607_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03608_ ) );
NAND3_X1 _10866_ ( .A1(_03603_ ), .A2(_03604_ ), .A3(_03608_ ), .ZN(_03609_ ) );
BUF_X4 _10867_ ( .A(_00968_ ), .Z(_03610_ ) );
BUF_X4 _10868_ ( .A(_03610_ ), .Z(_03611_ ) );
BUF_X4 _10869_ ( .A(_03611_ ), .Z(_03612_ ) );
BUF_X4 _10870_ ( .A(_03612_ ), .Z(_03613_ ) );
AND2_X1 _10871_ ( .A1(_00928_ ), .A2(\u_idu.imm_auipc_lui [20] ), .ZN(_03614_ ) );
BUF_X4 _10872_ ( .A(_03614_ ), .Z(_03615_ ) );
BUF_X4 _10873_ ( .A(_03615_ ), .Z(_03616_ ) );
AOI22_X1 _10874_ ( .A1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03613_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03617_ ) );
AND3_X1 _10875_ ( .A1(_03605_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03618_ ) );
BUF_X4 _10876_ ( .A(_03532_ ), .Z(_03619_ ) );
BUF_X4 _10877_ ( .A(_03619_ ), .Z(_03620_ ) );
BUF_X4 _10878_ ( .A(_03620_ ), .Z(_03621_ ) );
AOI21_X1 _10879_ ( .A(_03618_ ), .B1(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03621_ ), .ZN(_03622_ ) );
BUF_X2 _10880_ ( .A(_03539_ ), .Z(_03623_ ) );
NAND3_X1 _10881_ ( .A1(_03617_ ), .A2(_03622_ ), .A3(_03623_ ), .ZN(_03624_ ) );
AND2_X1 _10882_ ( .A1(_03624_ ), .A2(_03538_ ), .ZN(_03625_ ) );
AOI21_X1 _10883_ ( .A(_03600_ ), .B1(_03609_ ), .B2(_03625_ ), .ZN(_03626_ ) );
OAI21_X1 _10884_ ( .A(_03516_ ), .B1(_03507_ ), .B2(_03626_ ), .ZN(_03627_ ) );
OR2_X2 _10885_ ( .A1(_03588_ ), .A2(_03627_ ), .ZN(_03628_ ) );
BUF_X4 _10886_ ( .A(_03500_ ), .Z(_03629_ ) );
AOI211_X1 _10887_ ( .A(_03586_ ), .B(_03587_ ), .C1(_03628_ ), .C2(_03629_ ), .ZN(_03630_ ) );
BUF_X4 _10888_ ( .A(_01493_ ), .Z(_03631_ ) );
NOR2_X1 _10889_ ( .A1(_01518_ ), .A2(_03631_ ), .ZN(_03632_ ) );
OAI21_X1 _10890_ ( .A(_00302_ ), .B1(_03630_ ), .B2(_03632_ ), .ZN(_03633_ ) );
NAND2_X1 _10891_ ( .A1(_03498_ ), .A2(_03633_ ), .ZN(_00162_ ) );
AND3_X1 _10892_ ( .A1(_01658_ ), .A2(_03580_ ), .A3(_01659_ ), .ZN(_03634_ ) );
NOR2_X1 _10893_ ( .A1(\ar_data [21] ), .A2(_03510_ ), .ZN(_03635_ ) );
AND3_X1 _10894_ ( .A1(_03548_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03636_ ) );
BUF_X4 _10895_ ( .A(_03610_ ), .Z(_03637_ ) );
AOI221_X4 _10896_ ( .A(_03636_ ), .B1(_03533_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03637_ ), .ZN(_03638_ ) );
NAND3_X1 _10897_ ( .A1(_03606_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03639_ ) );
NAND3_X1 _10898_ ( .A1(_03638_ ), .A2(_03556_ ), .A3(_03639_ ), .ZN(_03640_ ) );
BUF_X4 _10899_ ( .A(_00926_ ), .Z(_03641_ ) );
AOI22_X1 _10900_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03612_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03642_ ) );
BUF_X4 _10901_ ( .A(_00980_ ), .Z(_03643_ ) );
BUF_X4 _10902_ ( .A(_03643_ ), .Z(_03644_ ) );
AOI22_X1 _10903_ ( .A1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03644_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03645_ ) );
NAND3_X1 _10904_ ( .A1(_03642_ ), .A2(_03645_ ), .A3(_03519_ ), .ZN(_03646_ ) );
AND3_X1 _10905_ ( .A1(_03640_ ), .A2(_03641_ ), .A3(_03646_ ), .ZN(_03647_ ) );
AND3_X1 _10906_ ( .A1(_03548_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03648_ ) );
AOI221_X4 _10907_ ( .A(_03648_ ), .B1(_03533_ ), .B2(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03552_ ), .ZN(_03649_ ) );
NAND3_X1 _10908_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03650_ ) );
NAND3_X1 _10909_ ( .A1(_03649_ ), .A2(_03623_ ), .A3(_03650_ ), .ZN(_03651_ ) );
OR3_X1 _10910_ ( .A1(_00925_ ), .A2(_03561_ ), .A3(_01624_ ), .ZN(_03652_ ) );
AOI21_X1 _10911_ ( .A(_03556_ ), .B1(_03652_ ), .B2(_03567_ ), .ZN(_03653_ ) );
BUF_X4 _10912_ ( .A(_03590_ ), .Z(_03654_ ) );
BUF_X4 _10913_ ( .A(_03654_ ), .Z(_03655_ ) );
NAND3_X1 _10914_ ( .A1(_03655_ ), .A2(_03562_ ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03656_ ) );
NAND3_X1 _10915_ ( .A1(_03571_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03657_ ) );
NAND3_X1 _10916_ ( .A1(_03653_ ), .A2(_03656_ ), .A3(_03657_ ), .ZN(_03658_ ) );
AND2_X1 _10917_ ( .A1(_03651_ ), .A2(_03658_ ), .ZN(_03659_ ) );
BUF_X4 _10918_ ( .A(_03537_ ), .Z(_03660_ ) );
BUF_X4 _10919_ ( .A(_03660_ ), .Z(_03661_ ) );
AOI21_X1 _10920_ ( .A(_03647_ ), .B1(_03659_ ), .B2(_03661_ ), .ZN(_03662_ ) );
OAI21_X1 _10921_ ( .A(_03516_ ), .B1(_03507_ ), .B2(_03662_ ), .ZN(_03663_ ) );
OR2_X2 _10922_ ( .A1(_03635_ ), .A2(_03663_ ), .ZN(_03664_ ) );
AOI211_X1 _10923_ ( .A(_03586_ ), .B(_03634_ ), .C1(_03664_ ), .C2(_03629_ ), .ZN(_03665_ ) );
AND2_X1 _10924_ ( .A1(_01664_ ), .A2(_02568_ ), .ZN(_03666_ ) );
OAI21_X1 _10925_ ( .A(_00302_ ), .B1(_03665_ ), .B2(_03666_ ), .ZN(_03667_ ) );
NAND2_X1 _10926_ ( .A1(_03498_ ), .A2(_03667_ ), .ZN(_00163_ ) );
AND3_X1 _10927_ ( .A1(_01714_ ), .A2(_03580_ ), .A3(_01716_ ), .ZN(_03668_ ) );
BUF_X4 _10928_ ( .A(_03515_ ), .Z(_03669_ ) );
BUF_X4 _10929_ ( .A(_03669_ ), .Z(_03670_ ) );
BUF_X16 _10930_ ( .A(_03510_ ), .Z(_03671_ ) );
BUF_X4 _10931_ ( .A(_03613_ ), .Z(_03672_ ) );
BUF_X4 _10932_ ( .A(_03534_ ), .Z(_03673_ ) );
AOI22_X1 _10933_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03672_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03674_ ) );
BUF_X4 _10934_ ( .A(_03517_ ), .Z(_03675_ ) );
BUF_X4 _10935_ ( .A(_03675_ ), .Z(_03676_ ) );
BUF_X4 _10936_ ( .A(_03676_ ), .Z(_03677_ ) );
BUF_X4 _10937_ ( .A(_03677_ ), .Z(_03678_ ) );
NAND3_X1 _10938_ ( .A1(_03607_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03679_ ) );
BUF_X4 _10939_ ( .A(_03606_ ), .Z(_03680_ ) );
NAND3_X1 _10940_ ( .A1(_03680_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03681_ ) );
NAND4_X1 _10941_ ( .A1(_03674_ ), .A2(_03678_ ), .A3(_03679_ ), .A4(_03681_ ), .ZN(_03682_ ) );
AOI22_X1 _10942_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03672_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03683_ ) );
BUF_X4 _10943_ ( .A(_03644_ ), .Z(_03684_ ) );
AOI22_X1 _10944_ ( .A1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03685_ ) );
NAND3_X1 _10945_ ( .A1(_03683_ ), .A2(_03685_ ), .A3(_03557_ ), .ZN(_03686_ ) );
BUF_X4 _10946_ ( .A(_03641_ ), .Z(_03687_ ) );
NAND3_X1 _10947_ ( .A1(_03682_ ), .A2(_03686_ ), .A3(_03687_ ), .ZN(_03688_ ) );
AND3_X1 _10948_ ( .A1(_03606_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03689_ ) );
BUF_X4 _10949_ ( .A(_03621_ ), .Z(_03690_ ) );
AOI21_X1 _10950_ ( .A(_03689_ ), .B1(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03690_ ), .ZN(_03691_ ) );
BUF_X4 _10951_ ( .A(_03655_ ), .Z(_03692_ ) );
NAND3_X1 _10952_ ( .A1(_03692_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03693_ ) );
NAND3_X1 _10953_ ( .A1(_03692_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03694_ ) );
NAND4_X1 _10954_ ( .A1(_03691_ ), .A2(_03557_ ), .A3(_03693_ ), .A4(_03694_ ), .ZN(_03695_ ) );
OR3_X1 _10955_ ( .A1(_00925_ ), .A2(_03562_ ), .A3(_01695_ ), .ZN(_03696_ ) );
AOI21_X1 _10956_ ( .A(_03601_ ), .B1(_03696_ ), .B2(_03567_ ), .ZN(_03697_ ) );
NAND3_X1 _10957_ ( .A1(_03559_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03698_ ) );
NAND3_X1 _10958_ ( .A1(_03607_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03699_ ) );
NAND3_X1 _10959_ ( .A1(_03697_ ), .A2(_03698_ ), .A3(_03699_ ), .ZN(_03700_ ) );
NAND2_X1 _10960_ ( .A1(_03695_ ), .A2(_03700_ ), .ZN(_03701_ ) );
OAI21_X1 _10961_ ( .A(_03688_ ), .B1(_03701_ ), .B2(_03687_ ), .ZN(_03702_ ) );
AOI21_X1 _10962_ ( .A(_03670_ ), .B1(_03671_ ), .B2(_03702_ ), .ZN(_03703_ ) );
BUF_X4 _10963_ ( .A(_03510_ ), .Z(_03704_ ) );
OAI21_X2 _10964_ ( .A(_03703_ ), .B1(\ar_data [20] ), .B2(_03704_ ), .ZN(_03705_ ) );
AOI211_X1 _10965_ ( .A(_03586_ ), .B(_03668_ ), .C1(_03705_ ), .C2(_03629_ ), .ZN(_03706_ ) );
AND2_X1 _10966_ ( .A1(_01722_ ), .A2(_02568_ ), .ZN(_03707_ ) );
OAI21_X1 _10967_ ( .A(_00302_ ), .B1(_03706_ ), .B2(_03707_ ), .ZN(_03708_ ) );
NAND2_X1 _10968_ ( .A1(_03498_ ), .A2(_03708_ ), .ZN(_00164_ ) );
AND3_X1 _10969_ ( .A1(_01773_ ), .A2(_03579_ ), .A3(_01775_ ), .ZN(_03709_ ) );
BUF_X8 _10970_ ( .A(_03509_ ), .Z(_03710_ ) );
AOI22_X1 _10971_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03637_ ), .B1(_03615_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03711_ ) );
AND3_X1 _10972_ ( .A1(_03548_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03712_ ) );
AOI21_X1 _10973_ ( .A(_03712_ ), .B1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03620_ ), .ZN(_03713_ ) );
AOI21_X1 _10974_ ( .A(_03539_ ), .B1(_03711_ ), .B2(_03713_ ), .ZN(_03714_ ) );
AND3_X1 _10975_ ( .A1(_03548_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03715_ ) );
AOI21_X1 _10976_ ( .A(_03715_ ), .B1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03637_ ), .ZN(_03716_ ) );
AOI22_X1 _10977_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03552_ ), .B1(_03533_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03717_ ) );
AOI21_X1 _10978_ ( .A(_03518_ ), .B1(_03716_ ), .B2(_03717_ ), .ZN(_03718_ ) );
OAI21_X1 _10979_ ( .A(_03641_ ), .B1(_03714_ ), .B2(_03718_ ), .ZN(_03719_ ) );
AND2_X1 _10980_ ( .A1(_00989_ ), .A2(fanout_net_20 ), .ZN(_03720_ ) );
BUF_X4 _10981_ ( .A(_03720_ ), .Z(_03721_ ) );
BUF_X4 _10982_ ( .A(_03721_ ), .Z(_03722_ ) );
AOI22_X1 _10983_ ( .A1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03644_ ), .B1(_03722_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03723_ ) );
AOI21_X1 _10984_ ( .A(_03518_ ), .B1(_03620_ ), .B2(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03724_ ) );
NAND3_X1 _10985_ ( .A1(_03654_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03725_ ) );
AND3_X1 _10986_ ( .A1(_03723_ ), .A2(_03724_ ), .A3(_03725_ ), .ZN(_03726_ ) );
AND3_X1 _10987_ ( .A1(_03590_ ), .A2(_03560_ ), .A3(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03727_ ) );
AOI21_X1 _10988_ ( .A(_03727_ ), .B1(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03722_ ), .ZN(_03728_ ) );
BUF_X4 _10989_ ( .A(_03521_ ), .Z(_03729_ ) );
AND2_X1 _10990_ ( .A1(_03549_ ), .A2(\u_reg.rf[1][19] ), .ZN(_03730_ ) );
OAI211_X1 _10991_ ( .A(_03728_ ), .B(_03676_ ), .C1(_03729_ ), .C2(_03730_ ), .ZN(_03731_ ) );
NAND2_X1 _10992_ ( .A1(_03731_ ), .A2(_03660_ ), .ZN(_03732_ ) );
OAI21_X1 _10993_ ( .A(_03719_ ), .B1(_03726_ ), .B2(_03732_ ), .ZN(_03733_ ) );
AOI21_X2 _10994_ ( .A(_03669_ ), .B1(_03710_ ), .B2(_03733_ ), .ZN(_03734_ ) );
OAI21_X2 _10995_ ( .A(_03734_ ), .B1(\ar_data [19] ), .B2(_03710_ ), .ZN(_03735_ ) );
AOI21_X1 _10996_ ( .A(_03709_ ), .B1(_03735_ ), .B2(_03500_ ), .ZN(_03736_ ) );
AOI22_X1 _10997_ ( .A1(_03736_ ), .A2(_03578_ ), .B1(_02362_ ), .B2(_01787_ ), .ZN(_03737_ ) );
NAND2_X4 _10998_ ( .A1(_03492_ ), .A2(_01505_ ), .ZN(_03738_ ) );
BUF_X4 _10999_ ( .A(_01106_ ), .Z(_03739_ ) );
BUF_X2 _11000_ ( .A(_01109_ ), .Z(_03740_ ) );
AOI22_X1 _11001_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_01787_ ), .ZN(_03741_ ) );
AOI221_X1 _11002_ ( .A(_02275_ ), .B1(_01090_ ), .B2(_03737_ ), .C1(_03738_ ), .C2(_03741_ ), .ZN(_00165_ ) );
AND3_X1 _11003_ ( .A1(_01840_ ), .A2(_03579_ ), .A3(_01841_ ), .ZN(_03742_ ) );
AOI22_X1 _11004_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03643_ ), .B1(_03532_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03743_ ) );
NAND3_X1 _11005_ ( .A1(_03520_ ), .A2(_03560_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03744_ ) );
NAND3_X1 _11006_ ( .A1(_03520_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03745_ ) );
AND4_X1 _11007_ ( .A1(_03675_ ), .A2(_03743_ ), .A3(_03744_ ), .A4(_03745_ ), .ZN(_03746_ ) );
NAND3_X1 _11008_ ( .A1(_03520_ ), .A2(_03560_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03747_ ) );
NAND3_X1 _11009_ ( .A1(_03527_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03748_ ) );
NAND3_X1 _11010_ ( .A1(_03527_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03749_ ) );
NAND3_X1 _11011_ ( .A1(_03747_ ), .A2(_03748_ ), .A3(_03749_ ), .ZN(_03750_ ) );
AOI211_X1 _11012_ ( .A(_03517_ ), .B(_03750_ ), .C1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03533_ ), .ZN(_03751_ ) );
OR3_X1 _11013_ ( .A1(_03746_ ), .A2(_03751_ ), .A3(_01028_ ), .ZN(_03752_ ) );
CLKBUF_X2 _11014_ ( .A(_00989_ ), .Z(_03753_ ) );
AND3_X1 _11015_ ( .A1(_03753_ ), .A2(_00978_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03754_ ) );
AOI221_X4 _11016_ ( .A(_03754_ ), .B1(_03532_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_03721_ ), .ZN(_03755_ ) );
NAND3_X1 _11017_ ( .A1(_03654_ ), .A2(_03561_ ), .A3(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03756_ ) );
AND3_X1 _11018_ ( .A1(_03755_ ), .A2(_03539_ ), .A3(_03756_ ), .ZN(_03757_ ) );
AOI22_X1 _11019_ ( .A1(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03637_ ), .B1(_03721_ ), .B2(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03758_ ) );
OAI21_X1 _11020_ ( .A(_00956_ ), .B1(_00958_ ), .B2(_01817_ ), .ZN(_03759_ ) );
NAND3_X1 _11021_ ( .A1(_03758_ ), .A2(_03676_ ), .A3(_03759_ ), .ZN(_03760_ ) );
NAND2_X1 _11022_ ( .A1(_03760_ ), .A2(_03537_ ), .ZN(_03761_ ) );
OAI21_X1 _11023_ ( .A(_03752_ ), .B1(_03757_ ), .B2(_03761_ ), .ZN(_03762_ ) );
AOI21_X1 _11024_ ( .A(_03515_ ), .B1(_03509_ ), .B2(_03762_ ), .ZN(_03763_ ) );
OAI21_X1 _11025_ ( .A(_03763_ ), .B1(\ar_data [18] ), .B2(_03710_ ), .ZN(_03764_ ) );
AOI211_X1 _11026_ ( .A(_03585_ ), .B(_03742_ ), .C1(_03764_ ), .C2(_03499_ ), .ZN(_03765_ ) );
AOI21_X1 _11027_ ( .A(_03765_ ), .B1(_02362_ ), .B2(_01852_ ), .ZN(_03766_ ) );
AOI22_X1 _11028_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_01852_ ), .ZN(_03767_ ) );
AOI221_X1 _11029_ ( .A(_02275_ ), .B1(_01090_ ), .B2(_03766_ ), .C1(_03738_ ), .C2(_03767_ ), .ZN(_00166_ ) );
NOR2_X2 _11030_ ( .A1(\ar_data [17] ), .A2(_03509_ ), .ZN(_03768_ ) );
AND3_X1 _11031_ ( .A1(_03528_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03769_ ) );
AOI21_X1 _11032_ ( .A(_03769_ ), .B1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03620_ ), .ZN(_03770_ ) );
NAND3_X1 _11033_ ( .A1(_03654_ ), .A2(_03561_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03771_ ) );
NAND3_X1 _11034_ ( .A1(_03605_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03772_ ) );
NAND4_X1 _11035_ ( .A1(_03770_ ), .A2(_03539_ ), .A3(_03771_ ), .A4(_03772_ ), .ZN(_03773_ ) );
AND3_X1 _11036_ ( .A1(_03527_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03774_ ) );
AOI21_X1 _11037_ ( .A(_03774_ ), .B1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03611_ ), .ZN(_03775_ ) );
AND2_X1 _11038_ ( .A1(_03548_ ), .A2(\u_reg.rf[1][17] ), .ZN(_03776_ ) );
OAI211_X1 _11039_ ( .A(_03775_ ), .B(_03675_ ), .C1(_03521_ ), .C2(_03776_ ), .ZN(_03777_ ) );
AND2_X1 _11040_ ( .A1(_03777_ ), .A2(_03537_ ), .ZN(_03778_ ) );
AOI21_X1 _11041_ ( .A(_03675_ ), .B1(_03620_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03779_ ) );
NAND3_X1 _11042_ ( .A1(_03605_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03780_ ) );
NAND3_X1 _11043_ ( .A1(_03654_ ), .A2(_03561_ ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03781_ ) );
NAND3_X1 _11044_ ( .A1(_03549_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03782_ ) );
NAND4_X1 _11045_ ( .A1(_03779_ ), .A2(_03780_ ), .A3(_03781_ ), .A4(_03782_ ), .ZN(_03783_ ) );
AND3_X1 _11046_ ( .A1(_00928_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03784_ ) );
AOI221_X4 _11047_ ( .A(_03784_ ), .B1(_00980_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03610_ ), .ZN(_03785_ ) );
AOI21_X1 _11048_ ( .A(_03555_ ), .B1(_03620_ ), .B2(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03786_ ) );
AOI21_X1 _11049_ ( .A(_03537_ ), .B1(_03785_ ), .B2(_03786_ ), .ZN(_03787_ ) );
AOI22_X1 _11050_ ( .A1(_03773_ ), .A2(_03778_ ), .B1(_03783_ ), .B2(_03787_ ), .ZN(_03788_ ) );
OAI21_X1 _11051_ ( .A(_03516_ ), .B1(_03507_ ), .B2(_03788_ ), .ZN(_03789_ ) );
OAI21_X1 _11052_ ( .A(_03499_ ), .B1(_03768_ ), .B2(_03789_ ), .ZN(_03790_ ) );
NAND3_X1 _11053_ ( .A1(_01896_ ), .A2(_03579_ ), .A3(_01897_ ), .ZN(_03791_ ) );
AND2_X1 _11054_ ( .A1(_03790_ ), .A2(_03791_ ), .ZN(_03792_ ) );
AOI22_X1 _11055_ ( .A1(_03792_ ), .A2(_03578_ ), .B1(_02362_ ), .B2(_01904_ ), .ZN(_03793_ ) );
AOI22_X1 _11056_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_01904_ ), .ZN(_03794_ ) );
AOI221_X1 _11057_ ( .A(_02454_ ), .B1(_01090_ ), .B2(_03793_ ), .C1(_03738_ ), .C2(_03794_ ), .ZN(_00167_ ) );
AND3_X1 _11058_ ( .A1(_01948_ ), .A2(_03579_ ), .A3(_01949_ ), .ZN(_03795_ ) );
AOI22_X1 _11059_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03637_ ), .B1(_03615_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03796_ ) );
AND3_X1 _11060_ ( .A1(_03548_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03797_ ) );
AOI21_X1 _11061_ ( .A(_03797_ ), .B1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03620_ ), .ZN(_03798_ ) );
AOI21_X1 _11062_ ( .A(_03676_ ), .B1(_03796_ ), .B2(_03798_ ), .ZN(_03799_ ) );
AOI22_X1 _11063_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03637_ ), .B1(_03615_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03800_ ) );
AOI22_X1 _11064_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03552_ ), .B1(_03533_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03801_ ) );
AOI21_X1 _11065_ ( .A(_03555_ ), .B1(_03800_ ), .B2(_03801_ ), .ZN(_03802_ ) );
OAI21_X1 _11066_ ( .A(_03641_ ), .B1(_03799_ ), .B2(_03802_ ), .ZN(_03803_ ) );
AOI22_X1 _11067_ ( .A1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03644_ ), .B1(_03722_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03804_ ) );
AOI21_X1 _11068_ ( .A(_03518_ ), .B1(_03620_ ), .B2(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03805_ ) );
NAND3_X1 _11069_ ( .A1(_03654_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03806_ ) );
AND3_X1 _11070_ ( .A1(_03804_ ), .A2(_03805_ ), .A3(_03806_ ), .ZN(_03807_ ) );
AND3_X1 _11071_ ( .A1(_03590_ ), .A2(_03560_ ), .A3(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03808_ ) );
AOI21_X1 _11072_ ( .A(_03808_ ), .B1(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03722_ ), .ZN(_03809_ ) );
AOI211_X1 _11073_ ( .A(_03523_ ), .B(_01929_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_03810_ ) );
OAI211_X1 _11074_ ( .A(_03809_ ), .B(_03676_ ), .C1(_03729_ ), .C2(_03810_ ), .ZN(_03811_ ) );
NAND2_X1 _11075_ ( .A1(_03811_ ), .A2(_03537_ ), .ZN(_03812_ ) );
OAI21_X1 _11076_ ( .A(_03803_ ), .B1(_03807_ ), .B2(_03812_ ), .ZN(_03813_ ) );
AOI21_X1 _11077_ ( .A(_03669_ ), .B1(_03509_ ), .B2(_03813_ ), .ZN(_03814_ ) );
OAI21_X2 _11078_ ( .A(_03814_ ), .B1(\ar_data [16] ), .B2(_03710_ ), .ZN(_03815_ ) );
AOI21_X1 _11079_ ( .A(_03795_ ), .B1(_03815_ ), .B2(_03500_ ), .ZN(_03816_ ) );
AOI22_X1 _11080_ ( .A1(_03816_ ), .A2(_03578_ ), .B1(_01490_ ), .B2(_01954_ ), .ZN(_03817_ ) );
AOI22_X1 _11081_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_01954_ ), .ZN(_03818_ ) );
AOI221_X1 _11082_ ( .A(_02454_ ), .B1(_01090_ ), .B2(_03817_ ), .C1(_03738_ ), .C2(_03818_ ), .ZN(_00168_ ) );
AND3_X1 _11083_ ( .A1(_01986_ ), .A2(_03579_ ), .A3(_01987_ ), .ZN(_03819_ ) );
AND3_X1 _11084_ ( .A1(_00957_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03820_ ) );
AOI221_X4 _11085_ ( .A(_03820_ ), .B1(_01019_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00968_ ), .ZN(_03821_ ) );
AOI21_X1 _11086_ ( .A(_00955_ ), .B1(_00980_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03822_ ) );
AOI21_X1 _11087_ ( .A(_01049_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03823_ ) );
AND3_X1 _11088_ ( .A1(_00957_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03824_ ) );
AOI221_X4 _11089_ ( .A(_03824_ ), .B1(_00980_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03610_ ), .ZN(_03825_ ) );
AOI221_X4 _11090_ ( .A(_01028_ ), .B1(_03821_ ), .B2(_03822_ ), .C1(_03823_ ), .C2(_03825_ ), .ZN(_03826_ ) );
AND3_X1 _11091_ ( .A1(_03753_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03827_ ) );
AOI21_X1 _11092_ ( .A(_03827_ ), .B1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03611_ ), .ZN(_03828_ ) );
AOI211_X1 _11093_ ( .A(_03560_ ), .B(_01968_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_03829_ ) );
OAI211_X1 _11094_ ( .A(_03828_ ), .B(_03675_ ), .C1(_03521_ ), .C2(_03829_ ), .ZN(_03830_ ) );
AOI22_X1 _11095_ ( .A1(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03643_ ), .B1(_03721_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03831_ ) );
AOI21_X1 _11096_ ( .A(_03517_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03832_ ) );
NAND3_X1 _11097_ ( .A1(_03590_ ), .A2(_03523_ ), .A3(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03833_ ) );
NAND3_X1 _11098_ ( .A1(_03831_ ), .A2(_03832_ ), .A3(_03833_ ), .ZN(_03834_ ) );
AND3_X1 _11099_ ( .A1(_03830_ ), .A2(_01028_ ), .A3(_03834_ ), .ZN(_03835_ ) );
OR2_X1 _11100_ ( .A1(_03826_ ), .A2(_03835_ ), .ZN(_03836_ ) );
AOI21_X1 _11101_ ( .A(_03515_ ), .B1(_03509_ ), .B2(_03836_ ), .ZN(_03837_ ) );
OAI21_X2 _11102_ ( .A(_03837_ ), .B1(\ar_data [15] ), .B2(_03710_ ), .ZN(_03838_ ) );
AOI211_X1 _11103_ ( .A(_03585_ ), .B(_03819_ ), .C1(_03838_ ), .C2(_03499_ ), .ZN(_03839_ ) );
AOI21_X1 _11104_ ( .A(_03839_ ), .B1(_02362_ ), .B2(_01994_ ), .ZN(_03840_ ) );
AOI22_X1 _11105_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_01994_ ), .ZN(_03841_ ) );
AOI221_X1 _11106_ ( .A(_02454_ ), .B1(_01090_ ), .B2(_03840_ ), .C1(_03738_ ), .C2(_03841_ ), .ZN(_00169_ ) );
AND3_X1 _11107_ ( .A1(_02042_ ), .A2(_03579_ ), .A3(_02043_ ), .ZN(_03842_ ) );
AOI22_X1 _11108_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03610_ ), .B1(_03615_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03843_ ) );
AND3_X1 _11109_ ( .A1(_03753_ ), .A2(_00978_ ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03844_ ) );
AOI21_X1 _11110_ ( .A(_03844_ ), .B1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03532_ ), .ZN(_03845_ ) );
AND3_X1 _11111_ ( .A1(_03843_ ), .A2(_03845_ ), .A3(_01049_ ), .ZN(_03846_ ) );
AOI21_X1 _11112_ ( .A(_03555_ ), .B1(_03620_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03847_ ) );
AND3_X1 _11113_ ( .A1(_03753_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03848_ ) );
AOI221_X4 _11114_ ( .A(_03848_ ), .B1(_00980_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03610_ ), .ZN(_03849_ ) );
AOI211_X1 _11115_ ( .A(_03537_ ), .B(_03846_ ), .C1(_03847_ ), .C2(_03849_ ), .ZN(_03850_ ) );
AOI22_X1 _11116_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03552_ ), .B1(_03721_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03851_ ) );
AOI21_X1 _11117_ ( .A(_03517_ ), .B1(_03533_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03852_ ) );
NAND3_X1 _11118_ ( .A1(_03590_ ), .A2(_03523_ ), .A3(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03853_ ) );
NAND3_X1 _11119_ ( .A1(_03851_ ), .A2(_03852_ ), .A3(_03853_ ), .ZN(_03854_ ) );
AOI22_X1 _11120_ ( .A1(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03611_ ), .B1(_03721_ ), .B2(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03855_ ) );
OAI21_X1 _11121_ ( .A(_00956_ ), .B1(_00958_ ), .B2(_02023_ ), .ZN(_03856_ ) );
NAND3_X1 _11122_ ( .A1(_03855_ ), .A2(_03675_ ), .A3(_03856_ ), .ZN(_03857_ ) );
AND3_X1 _11123_ ( .A1(_03854_ ), .A2(_03857_ ), .A3(_03537_ ), .ZN(_03858_ ) );
OR2_X1 _11124_ ( .A1(_03850_ ), .A2(_03858_ ), .ZN(_03859_ ) );
AOI21_X1 _11125_ ( .A(_03669_ ), .B1(_03509_ ), .B2(_03859_ ), .ZN(_03860_ ) );
OAI21_X2 _11126_ ( .A(_03860_ ), .B1(\ar_data [14] ), .B2(_03710_ ), .ZN(_03861_ ) );
AOI21_X1 _11127_ ( .A(_03842_ ), .B1(_03861_ ), .B2(_03500_ ), .ZN(_03862_ ) );
AOI22_X1 _11128_ ( .A1(_03862_ ), .A2(_03578_ ), .B1(_01490_ ), .B2(_02050_ ), .ZN(_03863_ ) );
AOI22_X1 _11129_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_02050_ ), .ZN(_03864_ ) );
AOI221_X1 _11130_ ( .A(_02454_ ), .B1(_01090_ ), .B2(_03863_ ), .C1(_03738_ ), .C2(_03864_ ), .ZN(_00170_ ) );
AND3_X1 _11131_ ( .A1(_02089_ ), .A2(_01440_ ), .A3(_02090_ ), .ZN(_03865_ ) );
AND3_X1 _11132_ ( .A1(_00989_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03866_ ) );
AOI221_X4 _11133_ ( .A(_03866_ ), .B1(_03532_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_00980_ ), .ZN(_03867_ ) );
NAND3_X1 _11134_ ( .A1(_03590_ ), .A2(_03523_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03868_ ) );
NAND3_X1 _11135_ ( .A1(_03867_ ), .A2(_03555_ ), .A3(_03868_ ), .ZN(_03869_ ) );
AND3_X1 _11136_ ( .A1(_03753_ ), .A2(fanout_net_20 ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03870_ ) );
AOI21_X1 _11137_ ( .A(_03870_ ), .B1(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03611_ ), .ZN(_03871_ ) );
AOI211_X1 _11138_ ( .A(_03560_ ), .B(_02070_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_03872_ ) );
OAI211_X1 _11139_ ( .A(_03871_ ), .B(_03675_ ), .C1(_03521_ ), .C2(_03872_ ), .ZN(_03873_ ) );
AND3_X1 _11140_ ( .A1(_03869_ ), .A2(_01028_ ), .A3(_03873_ ), .ZN(_03874_ ) );
NAND3_X1 _11141_ ( .A1(_03753_ ), .A2(_00978_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03875_ ) );
NAND3_X1 _11142_ ( .A1(_00928_ ), .A2(_00749_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03876_ ) );
NAND3_X1 _11143_ ( .A1(_00989_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03877_ ) );
AND3_X1 _11144_ ( .A1(_03875_ ), .A2(_03876_ ), .A3(_03877_ ), .ZN(_03878_ ) );
AOI21_X1 _11145_ ( .A(_01049_ ), .B1(_03532_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03879_ ) );
AOI21_X1 _11146_ ( .A(_03517_ ), .B1(_03532_ ), .B2(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03880_ ) );
NAND3_X1 _11147_ ( .A1(_03520_ ), .A2(_00749_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03881_ ) );
NAND3_X1 _11148_ ( .A1(_00928_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03882_ ) );
NAND3_X1 _11149_ ( .A1(_03753_ ), .A2(_00978_ ), .A3(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03883_ ) );
AND3_X1 _11150_ ( .A1(_03881_ ), .A2(_03882_ ), .A3(_03883_ ), .ZN(_03884_ ) );
AOI221_X4 _11151_ ( .A(_01028_ ), .B1(_03878_ ), .B2(_03879_ ), .C1(_03880_ ), .C2(_03884_ ), .ZN(_03885_ ) );
OR2_X1 _11152_ ( .A1(_03874_ ), .A2(_03885_ ), .ZN(_03886_ ) );
AOI21_X1 _11153_ ( .A(_03515_ ), .B1(_03509_ ), .B2(_03886_ ), .ZN(_03887_ ) );
OAI21_X2 _11154_ ( .A(_03887_ ), .B1(\ar_data [13] ), .B2(_03710_ ), .ZN(_03888_ ) );
AOI211_X1 _11155_ ( .A(_03585_ ), .B(_03865_ ), .C1(_03888_ ), .C2(_03499_ ), .ZN(_03889_ ) );
AOI21_X1 _11156_ ( .A(_03889_ ), .B1(_02362_ ), .B2(_02097_ ), .ZN(_03890_ ) );
AOI22_X1 _11157_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_02097_ ), .ZN(_03891_ ) );
AOI221_X1 _11158_ ( .A(_02454_ ), .B1(_01055_ ), .B2(_03890_ ), .C1(_03738_ ), .C2(_03891_ ), .ZN(_00171_ ) );
AND3_X1 _11159_ ( .A1(_02131_ ), .A2(_03579_ ), .A3(_02136_ ), .ZN(_03892_ ) );
AND3_X1 _11160_ ( .A1(_00957_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03893_ ) );
AOI221_X4 _11161_ ( .A(_03893_ ), .B1(_01019_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03610_ ), .ZN(_03894_ ) );
AOI21_X1 _11162_ ( .A(_03517_ ), .B1(_03643_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03895_ ) );
AOI21_X1 _11163_ ( .A(_01049_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03896_ ) );
AOI22_X1 _11164_ ( .A1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_00980_ ), .B1(_03610_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03897_ ) );
NAND3_X1 _11165_ ( .A1(_03527_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03898_ ) );
AND2_X1 _11166_ ( .A1(_03897_ ), .A2(_03898_ ), .ZN(_03899_ ) );
AOI221_X4 _11167_ ( .A(_01028_ ), .B1(_03894_ ), .B2(_03895_ ), .C1(_03896_ ), .C2(_03899_ ), .ZN(_03900_ ) );
AND3_X1 _11168_ ( .A1(_03753_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03901_ ) );
AOI21_X1 _11169_ ( .A(_03901_ ), .B1(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03611_ ), .ZN(_03902_ ) );
AND2_X1 _11170_ ( .A1(_03548_ ), .A2(\u_reg.rf[1][12] ), .ZN(_03903_ ) );
OAI211_X1 _11171_ ( .A(_03902_ ), .B(_03675_ ), .C1(_03521_ ), .C2(_03903_ ), .ZN(_03904_ ) );
AOI21_X1 _11172_ ( .A(_03517_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03905_ ) );
NAND3_X1 _11173_ ( .A1(_03590_ ), .A2(_03523_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03906_ ) );
NAND3_X1 _11174_ ( .A1(_03528_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03907_ ) );
NAND3_X1 _11175_ ( .A1(_03528_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03908_ ) );
NAND4_X1 _11176_ ( .A1(_03905_ ), .A2(_03906_ ), .A3(_03907_ ), .A4(_03908_ ), .ZN(_03909_ ) );
AND3_X1 _11177_ ( .A1(_03904_ ), .A2(_03909_ ), .A3(_01028_ ), .ZN(_03910_ ) );
OR2_X1 _11178_ ( .A1(_03900_ ), .A2(_03910_ ), .ZN(_03911_ ) );
AOI21_X1 _11179_ ( .A(_03515_ ), .B1(_03509_ ), .B2(_03911_ ), .ZN(_03912_ ) );
AND2_X1 _11180_ ( .A1(_02108_ ), .A2(_02110_ ), .ZN(\ar_data [12] ) );
OAI21_X2 _11181_ ( .A(_03912_ ), .B1(\ar_data [12] ), .B2(_03710_ ), .ZN(_03913_ ) );
AOI21_X1 _11182_ ( .A(_03892_ ), .B1(_03913_ ), .B2(_03500_ ), .ZN(_03914_ ) );
AOI22_X1 _11183_ ( .A1(_03914_ ), .A2(_03578_ ), .B1(_01490_ ), .B2(_02141_ ), .ZN(_03915_ ) );
AOI22_X1 _11184_ ( .A1(_03739_ ), .A2(_03740_ ), .B1(_03493_ ), .B2(_02141_ ), .ZN(_03916_ ) );
AOI221_X1 _11185_ ( .A(_02454_ ), .B1(_01055_ ), .B2(_03915_ ), .C1(_03738_ ), .C2(_03916_ ), .ZN(_00172_ ) );
AND3_X1 _11186_ ( .A1(_02171_ ), .A2(_03580_ ), .A3(_02172_ ), .ZN(_03917_ ) );
AOI22_X1 _11187_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03553_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03918_ ) );
AOI21_X1 _11188_ ( .A(_03539_ ), .B1(_03534_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03919_ ) );
NAND3_X1 _11189_ ( .A1(_03606_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03920_ ) );
AND3_X1 _11190_ ( .A1(_03918_ ), .A2(_03919_ ), .A3(_03920_ ), .ZN(_03921_ ) );
NAND3_X1 _11191_ ( .A1(_03529_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03922_ ) );
NAND2_X1 _11192_ ( .A1(_03922_ ), .A2(_03539_ ), .ZN(_03923_ ) );
NAND3_X1 _11193_ ( .A1(_03522_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03924_ ) );
NAND3_X1 _11194_ ( .A1(_03522_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03925_ ) );
NAND2_X1 _11195_ ( .A1(_03924_ ), .A2(_03925_ ), .ZN(_03926_ ) );
AOI211_X1 _11196_ ( .A(_03923_ ), .B(_03926_ ), .C1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03535_ ), .ZN(_03927_ ) );
OR3_X1 _11197_ ( .A1(_03921_ ), .A2(_03927_ ), .A3(_03538_ ), .ZN(_03928_ ) );
BUF_X4 _11198_ ( .A(_03722_ ), .Z(_03929_ ) );
AOI22_X1 _11199_ ( .A1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03929_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03930_ ) );
AOI21_X1 _11200_ ( .A(_03677_ ), .B1(_03690_ ), .B2(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03931_ ) );
NAND3_X1 _11201_ ( .A1(_03559_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03932_ ) );
AND3_X1 _11202_ ( .A1(_03930_ ), .A2(_03931_ ), .A3(_03932_ ), .ZN(_03933_ ) );
AND3_X1 _11203_ ( .A1(_03729_ ), .A2(_03543_ ), .A3(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03934_ ) );
AOI21_X1 _11204_ ( .A(_03934_ ), .B1(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03929_ ), .ZN(_03935_ ) );
AOI211_X1 _11205_ ( .A(_03569_ ), .B(_02152_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_03936_ ) );
OAI211_X1 _11206_ ( .A(_03935_ ), .B(_03678_ ), .C1(_03559_ ), .C2(_03936_ ), .ZN(_03937_ ) );
NAND2_X1 _11207_ ( .A1(_03937_ ), .A2(_03661_ ), .ZN(_03938_ ) );
OAI21_X1 _11208_ ( .A(_03928_ ), .B1(_03933_ ), .B2(_03938_ ), .ZN(_03939_ ) );
AOI21_X1 _11209_ ( .A(_03670_ ), .B1(_03671_ ), .B2(_03939_ ), .ZN(_03940_ ) );
OAI21_X1 _11210_ ( .A(_03940_ ), .B1(\ar_data [29] ), .B2(_03704_ ), .ZN(_03941_ ) );
AOI211_X1 _11211_ ( .A(_03586_ ), .B(_03917_ ), .C1(_03941_ ), .C2(_03629_ ), .ZN(_03942_ ) );
NOR2_X1 _11212_ ( .A1(_02177_ ), .A2(_03631_ ), .ZN(_03943_ ) );
OAI21_X1 _11213_ ( .A(_00302_ ), .B1(_03942_ ), .B2(_03943_ ), .ZN(_03944_ ) );
NAND2_X1 _11214_ ( .A1(_03498_ ), .A2(_03944_ ), .ZN(_00173_ ) );
BUF_X8 _11215_ ( .A(_03492_ ), .Z(_03945_ ) );
BUF_X4 _11216_ ( .A(_03493_ ), .Z(_03946_ ) );
OAI211_X1 _11217_ ( .A(_01070_ ), .B(_02227_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_03947_ ) );
AND3_X1 _11218_ ( .A1(_02211_ ), .A2(_03580_ ), .A3(_02217_ ), .ZN(_03948_ ) );
NAND3_X1 _11219_ ( .A1(_03522_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03949_ ) );
NAND3_X1 _11220_ ( .A1(_03529_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03950_ ) );
NAND2_X1 _11221_ ( .A1(_03949_ ), .A2(_03950_ ), .ZN(_03951_ ) );
AND3_X1 _11222_ ( .A1(_03528_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03952_ ) );
OR2_X1 _11223_ ( .A1(_03952_ ), .A2(_03518_ ), .ZN(_03953_ ) );
AOI211_X1 _11224_ ( .A(_03951_ ), .B(_03953_ ), .C1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03535_ ), .ZN(_03954_ ) );
AOI21_X1 _11225_ ( .A(_03601_ ), .B1(_03690_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03955_ ) );
AND3_X1 _11226_ ( .A1(_03549_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03956_ ) );
AOI221_X4 _11227_ ( .A(_03956_ ), .B1(_03644_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03612_ ), .ZN(_03957_ ) );
AOI211_X1 _11228_ ( .A(_03538_ ), .B(_03954_ ), .C1(_03955_ ), .C2(_03957_ ), .ZN(_03958_ ) );
OR3_X1 _11229_ ( .A1(_00925_ ), .A2(_03523_ ), .A3(_02196_ ), .ZN(_03959_ ) );
AOI21_X1 _11230_ ( .A(_03555_ ), .B1(_03959_ ), .B2(_00956_ ), .ZN(_03960_ ) );
AOI22_X1 _11231_ ( .A1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03612_ ), .B1(_03722_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03961_ ) );
AND3_X1 _11232_ ( .A1(_03527_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03962_ ) );
AOI221_X4 _11233_ ( .A(_03962_ ), .B1(_03643_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03637_ ), .ZN(_03963_ ) );
AOI21_X1 _11234_ ( .A(_03676_ ), .B1(_03534_ ), .B2(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03964_ ) );
AOI221_X4 _11235_ ( .A(_03641_ ), .B1(_03960_ ), .B2(_03961_ ), .C1(_03963_ ), .C2(_03964_ ), .ZN(_03965_ ) );
OR2_X1 _11236_ ( .A1(_03958_ ), .A2(_03965_ ), .ZN(_03966_ ) );
AOI21_X1 _11237_ ( .A(_03670_ ), .B1(_03671_ ), .B2(_03966_ ), .ZN(_03967_ ) );
OAI21_X1 _11238_ ( .A(_03967_ ), .B1(\ar_data [11] ), .B2(_03704_ ), .ZN(_03968_ ) );
AOI211_X1 _11239_ ( .A(_03586_ ), .B(_03948_ ), .C1(_03968_ ), .C2(_03629_ ), .ZN(_03969_ ) );
NOR2_X1 _11240_ ( .A1(_03631_ ), .A2(_02226_ ), .ZN(_03970_ ) );
OAI21_X1 _11241_ ( .A(_00302_ ), .B1(_03969_ ), .B2(_03970_ ), .ZN(_03971_ ) );
NAND2_X1 _11242_ ( .A1(_03947_ ), .A2(_03971_ ), .ZN(_00174_ ) );
OAI211_X1 _11243_ ( .A(_01069_ ), .B(_02273_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_03972_ ) );
BUF_X4 _11244_ ( .A(_03585_ ), .Z(_03973_ ) );
CLKBUF_X2 _11245_ ( .A(_03579_ ), .Z(_03974_ ) );
AND3_X1 _11246_ ( .A1(_02265_ ), .A2(_03974_ ), .A3(_02266_ ), .ZN(_03975_ ) );
AND3_X1 _11247_ ( .A1(_03520_ ), .A2(_00749_ ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03976_ ) );
AOI221_X4 _11248_ ( .A(_03976_ ), .B1(_03643_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_03615_ ), .ZN(_03977_ ) );
AOI21_X1 _11249_ ( .A(_03555_ ), .B1(_03620_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03978_ ) );
AOI21_X1 _11250_ ( .A(_03518_ ), .B1(_03534_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03979_ ) );
AND3_X1 _11251_ ( .A1(_03520_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03980_ ) );
AOI221_X4 _11252_ ( .A(_03980_ ), .B1(_03643_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03611_ ), .ZN(_03981_ ) );
AOI221_X4 _11253_ ( .A(_03537_ ), .B1(_03977_ ), .B2(_03978_ ), .C1(_03979_ ), .C2(_03981_ ), .ZN(_03982_ ) );
AND3_X1 _11254_ ( .A1(_03527_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03983_ ) );
AOI221_X4 _11255_ ( .A(_03983_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03552_ ), .ZN(_03984_ ) );
NAND3_X1 _11256_ ( .A1(_03655_ ), .A2(_03562_ ), .A3(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03985_ ) );
NAND3_X1 _11257_ ( .A1(_03984_ ), .A2(_03556_ ), .A3(_03985_ ), .ZN(_03986_ ) );
AOI22_X1 _11258_ ( .A1(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03612_ ), .B1(_03722_ ), .B2(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03987_ ) );
OAI21_X1 _11259_ ( .A(_00956_ ), .B1(_00958_ ), .B2(_02245_ ), .ZN(_03988_ ) );
NAND3_X1 _11260_ ( .A1(_03987_ ), .A2(_03519_ ), .A3(_03988_ ), .ZN(_03989_ ) );
AND3_X1 _11261_ ( .A1(_03986_ ), .A2(_03989_ ), .A3(_03660_ ), .ZN(_03990_ ) );
OR2_X1 _11262_ ( .A1(_03982_ ), .A2(_03990_ ), .ZN(_03991_ ) );
AOI21_X2 _11263_ ( .A(_03669_ ), .B1(_03511_ ), .B2(_03991_ ), .ZN(_03992_ ) );
AND2_X1 _11264_ ( .A1(_02236_ ), .A2(_02238_ ), .ZN(\ar_data [10] ) );
OAI21_X2 _11265_ ( .A(_03992_ ), .B1(\ar_data [10] ), .B2(_03671_ ), .ZN(_03993_ ) );
BUF_X4 _11266_ ( .A(_03500_ ), .Z(_03994_ ) );
AOI211_X1 _11267_ ( .A(_03973_ ), .B(_03975_ ), .C1(_03993_ ), .C2(_03994_ ), .ZN(_03995_ ) );
AOI21_X1 _11268_ ( .A(_03995_ ), .B1(_02568_ ), .B2(_02273_ ), .ZN(_03996_ ) );
OAI21_X1 _11269_ ( .A(_03972_ ), .B1(_01854_ ), .B2(_03996_ ), .ZN(_00175_ ) );
OAI211_X1 _11270_ ( .A(_01070_ ), .B(_02316_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_03997_ ) );
BUF_X4 _11271_ ( .A(_01569_ ), .Z(_03998_ ) );
AND3_X1 _11272_ ( .A1(_02311_ ), .A2(_03580_ ), .A3(_02312_ ), .ZN(_03999_ ) );
AND3_X1 _11273_ ( .A1(_03527_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04000_ ) );
AOI221_X4 _11274_ ( .A(_04000_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03611_ ), .ZN(_04001_ ) );
AOI21_X1 _11275_ ( .A(_03518_ ), .B1(_03644_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04002_ ) );
AOI21_X1 _11276_ ( .A(_03539_ ), .B1(_03621_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04003_ ) );
AOI22_X1 _11277_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03552_ ), .B1(_03637_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04004_ ) );
NAND3_X1 _11278_ ( .A1(_03605_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04005_ ) );
AND2_X1 _11279_ ( .A1(_04004_ ), .A2(_04005_ ), .ZN(_04006_ ) );
AOI221_X4 _11280_ ( .A(_03660_ ), .B1(_04001_ ), .B2(_04002_ ), .C1(_04003_ ), .C2(_04006_ ), .ZN(_04007_ ) );
AOI22_X1 _11281_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03553_ ), .B1(_03929_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04008_ ) );
AOI21_X1 _11282_ ( .A(_03676_ ), .B1(_03621_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04009_ ) );
NAND3_X1 _11283_ ( .A1(_03655_ ), .A2(_03562_ ), .A3(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04010_ ) );
NAND3_X1 _11284_ ( .A1(_04008_ ), .A2(_04009_ ), .A3(_04010_ ), .ZN(_04011_ ) );
AOI22_X1 _11285_ ( .A1(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03613_ ), .B1(_03929_ ), .B2(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04012_ ) );
OAI21_X1 _11286_ ( .A(_00956_ ), .B1(_00958_ ), .B2(_02293_ ), .ZN(_04013_ ) );
NAND3_X1 _11287_ ( .A1(_04012_ ), .A2(_03677_ ), .A3(_04013_ ), .ZN(_04014_ ) );
AND3_X1 _11288_ ( .A1(_04011_ ), .A2(_04014_ ), .A3(_03660_ ), .ZN(_04015_ ) );
OR2_X1 _11289_ ( .A1(_04007_ ), .A2(_04015_ ), .ZN(_04016_ ) );
AOI21_X1 _11290_ ( .A(_03670_ ), .B1(_03671_ ), .B2(_04016_ ), .ZN(_04017_ ) );
AND2_X1 _11291_ ( .A1(_02284_ ), .A2(_02286_ ), .ZN(\ar_data [9] ) );
OAI21_X2 _11292_ ( .A(_04017_ ), .B1(\ar_data [9] ), .B2(_03704_ ), .ZN(_04018_ ) );
AOI211_X1 _11293_ ( .A(_03586_ ), .B(_03999_ ), .C1(_04018_ ), .C2(_03629_ ), .ZN(_04019_ ) );
NOR3_X1 _11294_ ( .A1(_03631_ ), .A2(_02359_ ), .A3(_00881_ ), .ZN(_04020_ ) );
OAI21_X1 _11295_ ( .A(_03998_ ), .B1(_04019_ ), .B2(_04020_ ), .ZN(_04021_ ) );
NAND2_X1 _11296_ ( .A1(_03997_ ), .A2(_04021_ ), .ZN(_00176_ ) );
OAI211_X1 _11297_ ( .A(_01069_ ), .B(_02360_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_04022_ ) );
AND3_X1 _11298_ ( .A1(_02352_ ), .A2(_03974_ ), .A3(_02353_ ), .ZN(_04023_ ) );
AOI21_X1 _11299_ ( .A(_03518_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04024_ ) );
NAND3_X1 _11300_ ( .A1(_03522_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04025_ ) );
NAND3_X1 _11301_ ( .A1(_03529_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04026_ ) );
NAND3_X1 _11302_ ( .A1(_03529_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04027_ ) );
AND4_X1 _11303_ ( .A1(_04024_ ), .A2(_04025_ ), .A3(_04026_ ), .A4(_04027_ ), .ZN(_04028_ ) );
AOI21_X1 _11304_ ( .A(_03623_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04029_ ) );
AND3_X1 _11305_ ( .A1(_03528_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04030_ ) );
AOI221_X4 _11306_ ( .A(_04030_ ), .B1(_03644_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03612_ ), .ZN(_04031_ ) );
AOI211_X1 _11307_ ( .A(_03660_ ), .B(_04028_ ), .C1(_04029_ ), .C2(_04031_ ), .ZN(_04032_ ) );
AOI22_X1 _11308_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03613_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04033_ ) );
AND3_X1 _11309_ ( .A1(_03549_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04034_ ) );
AOI21_X1 _11310_ ( .A(_04034_ ), .B1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03534_ ), .ZN(_04035_ ) );
NAND3_X1 _11311_ ( .A1(_04033_ ), .A2(_04035_ ), .A3(_03556_ ), .ZN(_04036_ ) );
AOI22_X1 _11312_ ( .A1(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03612_ ), .B1(_03722_ ), .B2(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04037_ ) );
OAI21_X1 _11313_ ( .A(_00956_ ), .B1(_00958_ ), .B2(_02333_ ), .ZN(_04038_ ) );
NAND3_X1 _11314_ ( .A1(_04037_ ), .A2(_03519_ ), .A3(_04038_ ), .ZN(_04039_ ) );
AND3_X1 _11315_ ( .A1(_04036_ ), .A2(_04039_ ), .A3(_03660_ ), .ZN(_04040_ ) );
OR2_X1 _11316_ ( .A1(_04032_ ), .A2(_04040_ ), .ZN(_04041_ ) );
AOI21_X2 _11317_ ( .A(_03669_ ), .B1(_03511_ ), .B2(_04041_ ), .ZN(_04042_ ) );
OAI21_X1 _11318_ ( .A(_04042_ ), .B1(\ar_data [8] ), .B2(_03671_ ), .ZN(_04043_ ) );
AOI211_X1 _11319_ ( .A(_03973_ ), .B(_04023_ ), .C1(_04043_ ), .C2(_03994_ ), .ZN(_04044_ ) );
AOI21_X1 _11320_ ( .A(_04044_ ), .B1(_02568_ ), .B2(_02360_ ), .ZN(_04045_ ) );
OAI21_X1 _11321_ ( .A(_04022_ ), .B1(_01854_ ), .B2(_04045_ ), .ZN(_00177_ ) );
OAI211_X1 _11322_ ( .A(_01070_ ), .B(_02387_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_04046_ ) );
AND3_X1 _11323_ ( .A1(_02396_ ), .A2(_03580_ ), .A3(_02397_ ), .ZN(_04047_ ) );
AOI22_X1 _11324_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03672_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04048_ ) );
AND3_X1 _11325_ ( .A1(_03541_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04049_ ) );
AOI21_X1 _11326_ ( .A(_04049_ ), .B1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03673_ ), .ZN(_04050_ ) );
NAND3_X1 _11327_ ( .A1(_04048_ ), .A2(_04050_ ), .A3(_03557_ ), .ZN(_04051_ ) );
AOI22_X1 _11328_ ( .A1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03613_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04052_ ) );
AOI21_X1 _11329_ ( .A(_03623_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04053_ ) );
NAND3_X1 _11330_ ( .A1(_03607_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04054_ ) );
NAND3_X1 _11331_ ( .A1(_04052_ ), .A2(_04053_ ), .A3(_04054_ ), .ZN(_04055_ ) );
NAND3_X1 _11332_ ( .A1(_04051_ ), .A2(_04055_ ), .A3(_03687_ ), .ZN(_04056_ ) );
NAND3_X1 _11333_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04057_ ) );
NAND3_X1 _11334_ ( .A1(_03571_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04058_ ) );
NAND3_X1 _11335_ ( .A1(_03571_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04059_ ) );
NAND3_X1 _11336_ ( .A1(_04057_ ), .A2(_04058_ ), .A3(_04059_ ), .ZN(_04060_ ) );
AOI211_X1 _11337_ ( .A(_03678_ ), .B(_04060_ ), .C1(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03690_ ), .ZN(_04061_ ) );
OR3_X1 _11338_ ( .A1(_00925_ ), .A2(_03543_ ), .A3(_02372_ ), .ZN(_04062_ ) );
AOI21_X1 _11339_ ( .A(_03623_ ), .B1(_04062_ ), .B2(_03567_ ), .ZN(_04063_ ) );
NAND3_X1 _11340_ ( .A1(_03692_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04064_ ) );
NAND3_X1 _11341_ ( .A1(_03607_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04065_ ) );
NAND3_X1 _11342_ ( .A1(_04063_ ), .A2(_04064_ ), .A3(_04065_ ), .ZN(_04066_ ) );
NAND2_X1 _11343_ ( .A1(_04066_ ), .A2(_03661_ ), .ZN(_04067_ ) );
OAI21_X1 _11344_ ( .A(_04056_ ), .B1(_04061_ ), .B2(_04067_ ), .ZN(_04068_ ) );
AOI21_X2 _11345_ ( .A(_03670_ ), .B1(_03511_ ), .B2(_04068_ ), .ZN(_04069_ ) );
BUF_X2 _11346_ ( .A(_03510_ ), .Z(_04070_ ) );
OAI21_X1 _11347_ ( .A(_04069_ ), .B1(\ar_data [7] ), .B2(_04070_ ), .ZN(_04071_ ) );
AOI211_X1 _11348_ ( .A(_03586_ ), .B(_04047_ ), .C1(_04071_ ), .C2(_03629_ ), .ZN(_04072_ ) );
NOR3_X1 _11349_ ( .A1(_01493_ ), .A2(_02359_ ), .A3(_00886_ ), .ZN(_04073_ ) );
OAI21_X1 _11350_ ( .A(_03998_ ), .B1(_04072_ ), .B2(_04073_ ), .ZN(_04074_ ) );
NAND2_X1 _11351_ ( .A1(_04046_ ), .A2(_04074_ ), .ZN(_00178_ ) );
OAI211_X1 _11352_ ( .A(_01069_ ), .B(_02452_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_04075_ ) );
AND3_X1 _11353_ ( .A1(_02447_ ), .A2(_03974_ ), .A3(_02448_ ), .ZN(_04076_ ) );
AOI22_X1 _11354_ ( .A1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03621_ ), .B2(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04077_ ) );
NAND3_X1 _11355_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04078_ ) );
NAND3_X1 _11356_ ( .A1(_03558_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04079_ ) );
NAND4_X1 _11357_ ( .A1(_04077_ ), .A2(_03677_ ), .A3(_04078_ ), .A4(_04079_ ), .ZN(_04080_ ) );
NAND3_X1 _11358_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04081_ ) );
INV_X1 _11359_ ( .A(_03684_ ), .ZN(_04082_ ) );
INV_X1 _11360_ ( .A(_03616_ ), .ZN(_04083_ ) );
OAI221_X1 _11361_ ( .A(_04081_ ), .B1(_04082_ ), .B2(_02405_ ), .C1(_02409_ ), .C2(_04083_ ), .ZN(_04084_ ) );
INV_X1 _11362_ ( .A(_03621_ ), .ZN(_04085_ ) );
OAI21_X1 _11363_ ( .A(_03601_ ), .B1(_04085_ ), .B2(_02402_ ), .ZN(_04086_ ) );
OAI211_X1 _11364_ ( .A(_03641_ ), .B(_04080_ ), .C1(_04084_ ), .C2(_04086_ ), .ZN(_04087_ ) );
AND3_X1 _11365_ ( .A1(_03529_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04088_ ) );
AOI21_X1 _11366_ ( .A(_04088_ ), .B1(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03621_ ), .ZN(_04089_ ) );
NAND3_X1 _11367_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04090_ ) );
NAND3_X1 _11368_ ( .A1(_03571_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04091_ ) );
AND4_X1 _11369_ ( .A1(_03601_ ), .A2(_04089_ ), .A3(_04090_ ), .A4(_04091_ ), .ZN(_04092_ ) );
OAI211_X1 _11370_ ( .A(\u_idu.imm_auipc_lui [20] ), .B(\u_reg.rf[1][6] ), .C1(_02563_ ), .C2(_01078_ ), .ZN(_04093_ ) );
AOI21_X1 _11371_ ( .A(_03623_ ), .B1(_04093_ ), .B2(_03567_ ), .ZN(_04094_ ) );
BUF_X4 _11372_ ( .A(_03729_ ), .Z(_04095_ ) );
BUF_X4 _11373_ ( .A(_03562_ ), .Z(_04096_ ) );
NAND3_X1 _11374_ ( .A1(_04095_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04097_ ) );
NAND3_X1 _11375_ ( .A1(_03680_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04098_ ) );
NAND3_X1 _11376_ ( .A1(_04094_ ), .A2(_04097_ ), .A3(_04098_ ), .ZN(_04099_ ) );
NAND2_X1 _11377_ ( .A1(_04099_ ), .A2(_03661_ ), .ZN(_04100_ ) );
OAI21_X1 _11378_ ( .A(_04087_ ), .B1(_04092_ ), .B2(_04100_ ), .ZN(_04101_ ) );
AOI21_X2 _11379_ ( .A(_03669_ ), .B1(_03510_ ), .B2(_04101_ ), .ZN(_04102_ ) );
OAI21_X1 _11380_ ( .A(_04102_ ), .B1(\ar_data [6] ), .B2(_03671_ ), .ZN(_04103_ ) );
AOI211_X1 _11381_ ( .A(_03973_ ), .B(_04076_ ), .C1(_04103_ ), .C2(_03994_ ), .ZN(_04104_ ) );
AOI21_X1 _11382_ ( .A(_04104_ ), .B1(_02568_ ), .B2(_02452_ ), .ZN(_04105_ ) );
OAI21_X1 _11383_ ( .A(_04075_ ), .B1(_01854_ ), .B2(_04105_ ), .ZN(_00179_ ) );
OAI211_X1 _11384_ ( .A(_01070_ ), .B(_02457_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_04106_ ) );
NOR3_X1 _11385_ ( .A1(_02499_ ), .A2(_03500_ ), .A3(_02510_ ), .ZN(_04107_ ) );
AOI22_X1 _11386_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03672_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04108_ ) );
AND3_X1 _11387_ ( .A1(_03541_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04109_ ) );
AOI21_X1 _11388_ ( .A(_04109_ ), .B1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03673_ ), .ZN(_04110_ ) );
NAND3_X1 _11389_ ( .A1(_04108_ ), .A2(_04110_ ), .A3(_03557_ ), .ZN(_04111_ ) );
AOI22_X1 _11390_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03672_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04112_ ) );
AOI22_X1 _11391_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03535_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04113_ ) );
NAND3_X1 _11392_ ( .A1(_04112_ ), .A2(_04113_ ), .A3(_03678_ ), .ZN(_04114_ ) );
NAND3_X1 _11393_ ( .A1(_04111_ ), .A2(_04114_ ), .A3(_03687_ ), .ZN(_04115_ ) );
NAND3_X1 _11394_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04116_ ) );
NAND3_X1 _11395_ ( .A1(_03571_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04117_ ) );
NAND3_X1 _11396_ ( .A1(_03571_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04118_ ) );
NAND3_X1 _11397_ ( .A1(_04116_ ), .A2(_04117_ ), .A3(_04118_ ), .ZN(_04119_ ) );
AOI211_X1 _11398_ ( .A(_03678_ ), .B(_04119_ ), .C1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03690_ ), .ZN(_04120_ ) );
AOI22_X1 _11399_ ( .A1(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03672_ ), .B1(_03929_ ), .B2(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04121_ ) );
OAI21_X1 _11400_ ( .A(_03567_ ), .B1(_00958_ ), .B2(_02476_ ), .ZN(_04122_ ) );
NAND3_X1 _11401_ ( .A1(_04121_ ), .A2(_03678_ ), .A3(_04122_ ), .ZN(_04123_ ) );
NAND2_X1 _11402_ ( .A1(_04123_ ), .A2(_03661_ ), .ZN(_04124_ ) );
OAI21_X1 _11403_ ( .A(_04115_ ), .B1(_04120_ ), .B2(_04124_ ), .ZN(_04125_ ) );
AOI21_X2 _11404_ ( .A(_03670_ ), .B1(_03511_ ), .B2(_04125_ ), .ZN(_04126_ ) );
OAI21_X1 _11405_ ( .A(_04126_ ), .B1(\ar_data [5] ), .B2(_04070_ ), .ZN(_04127_ ) );
AOI211_X1 _11406_ ( .A(_03586_ ), .B(_04107_ ), .C1(_04127_ ), .C2(_03629_ ), .ZN(_04128_ ) );
NOR3_X1 _11407_ ( .A1(_01493_ ), .A2(_02359_ ), .A3(_00656_ ), .ZN(_04129_ ) );
OAI21_X1 _11408_ ( .A(_03998_ ), .B1(_04128_ ), .B2(_04129_ ), .ZN(_04130_ ) );
NAND2_X1 _11409_ ( .A1(_04106_ ), .A2(_04130_ ), .ZN(_00180_ ) );
OAI211_X1 _11410_ ( .A(_01070_ ), .B(_02566_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_04131_ ) );
AND3_X1 _11411_ ( .A1(_02556_ ), .A2(_03974_ ), .A3(_02557_ ), .ZN(_04132_ ) );
AND3_X1 _11412_ ( .A1(_03521_ ), .A2(_03561_ ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04133_ ) );
AOI221_X4 _11413_ ( .A(_04133_ ), .B1(_03722_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03644_ ), .ZN(_04134_ ) );
OAI211_X1 _11414_ ( .A(_04134_ ), .B(_03557_ ), .C1(_02537_ ), .C2(_04085_ ), .ZN(_04135_ ) );
AND3_X1 _11415_ ( .A1(_03605_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04136_ ) );
AND3_X1 _11416_ ( .A1(_03654_ ), .A2(_03561_ ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04137_ ) );
OR2_X1 _11417_ ( .A1(_04136_ ), .A2(_04137_ ), .ZN(_04138_ ) );
AOI21_X1 _11418_ ( .A(_03655_ ), .B1(\u_reg.rf[1][4] ), .B2(_03606_ ), .ZN(_04139_ ) );
OR3_X1 _11419_ ( .A1(_04138_ ), .A2(_03623_ ), .A3(_04139_ ), .ZN(_04140_ ) );
NAND3_X1 _11420_ ( .A1(_04135_ ), .A2(_03661_ ), .A3(_04140_ ), .ZN(_04141_ ) );
AOI22_X1 _11421_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03672_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04142_ ) );
AND3_X1 _11422_ ( .A1(_03606_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04143_ ) );
AOI21_X1 _11423_ ( .A(_04143_ ), .B1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03690_ ), .ZN(_04144_ ) );
NAND3_X1 _11424_ ( .A1(_04142_ ), .A2(_04144_ ), .A3(_03557_ ), .ZN(_04145_ ) );
AOI22_X1 _11425_ ( .A1(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03672_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04146_ ) );
AOI21_X1 _11426_ ( .A(_03623_ ), .B1(_03690_ ), .B2(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04147_ ) );
NAND3_X1 _11427_ ( .A1(_03607_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04148_ ) );
NAND3_X1 _11428_ ( .A1(_04146_ ), .A2(_04147_ ), .A3(_04148_ ), .ZN(_04149_ ) );
NAND3_X1 _11429_ ( .A1(_04145_ ), .A2(_04149_ ), .A3(_03687_ ), .ZN(_04150_ ) );
NAND2_X1 _11430_ ( .A1(_04141_ ), .A2(_04150_ ), .ZN(_04151_ ) );
AOI21_X2 _11431_ ( .A(_03669_ ), .B1(_03511_ ), .B2(_04151_ ), .ZN(_04152_ ) );
OAI21_X1 _11432_ ( .A(_04152_ ), .B1(\ar_data [4] ), .B2(_03704_ ), .ZN(_04153_ ) );
AOI211_X1 _11433_ ( .A(_03586_ ), .B(_04132_ ), .C1(_04153_ ), .C2(_03629_ ), .ZN(_04154_ ) );
AND2_X1 _11434_ ( .A1(_02568_ ), .A2(_02566_ ), .ZN(_04155_ ) );
OAI21_X1 _11435_ ( .A(_03998_ ), .B1(_04154_ ), .B2(_04155_ ), .ZN(_04156_ ) );
NAND2_X1 _11436_ ( .A1(_04131_ ), .A2(_04156_ ), .ZN(_00181_ ) );
OAI211_X1 _11437_ ( .A(_01069_ ), .B(_02616_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_04157_ ) );
AND3_X1 _11438_ ( .A1(_02609_ ), .A2(_03974_ ), .A3(_02610_ ), .ZN(_04158_ ) );
AOI22_X1 _11439_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03613_ ), .B1(_03616_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04159_ ) );
AND3_X1 _11440_ ( .A1(_03541_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04160_ ) );
AOI21_X1 _11441_ ( .A(_04160_ ), .B1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03535_ ), .ZN(_04161_ ) );
NAND3_X1 _11442_ ( .A1(_04159_ ), .A2(_04161_ ), .A3(_03601_ ), .ZN(_04162_ ) );
AOI22_X1 _11443_ ( .A1(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03613_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04163_ ) );
AOI21_X1 _11444_ ( .A(_03556_ ), .B1(_03535_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04164_ ) );
NAND3_X1 _11445_ ( .A1(_03680_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04165_ ) );
NAND3_X1 _11446_ ( .A1(_04163_ ), .A2(_04164_ ), .A3(_04165_ ), .ZN(_04166_ ) );
NAND3_X1 _11447_ ( .A1(_04162_ ), .A2(_04166_ ), .A3(_03641_ ), .ZN(_04167_ ) );
AOI21_X1 _11448_ ( .A(_03519_ ), .B1(_03535_ ), .B2(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04168_ ) );
NAND3_X1 _11449_ ( .A1(_04095_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04169_ ) );
NAND3_X1 _11450_ ( .A1(_03571_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04170_ ) );
NAND3_X1 _11451_ ( .A1(_03571_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04171_ ) );
AND4_X1 _11452_ ( .A1(_04168_ ), .A2(_04169_ ), .A3(_04170_ ), .A4(_04171_ ), .ZN(_04172_ ) );
OR3_X1 _11453_ ( .A1(_00925_ ), .A2(_03524_ ), .A3(_02586_ ), .ZN(_04173_ ) );
AOI21_X1 _11454_ ( .A(_03556_ ), .B1(_04173_ ), .B2(_03567_ ), .ZN(_04174_ ) );
NAND3_X1 _11455_ ( .A1(_04095_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04175_ ) );
NAND3_X1 _11456_ ( .A1(_03680_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04176_ ) );
NAND3_X1 _11457_ ( .A1(_04174_ ), .A2(_04175_ ), .A3(_04176_ ), .ZN(_04177_ ) );
NAND2_X1 _11458_ ( .A1(_04177_ ), .A2(_03661_ ), .ZN(_04178_ ) );
OAI21_X1 _11459_ ( .A(_04167_ ), .B1(_04172_ ), .B2(_04178_ ), .ZN(_04179_ ) );
AOI21_X2 _11460_ ( .A(_03669_ ), .B1(_03510_ ), .B2(_04179_ ), .ZN(_04180_ ) );
OAI21_X1 _11461_ ( .A(_04180_ ), .B1(\ar_data [3] ), .B2(_03671_ ), .ZN(_04181_ ) );
AOI211_X1 _11462_ ( .A(_03973_ ), .B(_04158_ ), .C1(_04181_ ), .C2(_03994_ ), .ZN(_04182_ ) );
AOI21_X1 _11463_ ( .A(_04182_ ), .B1(_02568_ ), .B2(_02616_ ), .ZN(_04183_ ) );
OAI21_X1 _11464_ ( .A(_04157_ ), .B1(_01854_ ), .B2(_04183_ ), .ZN(_00182_ ) );
AOI22_X1 _11465_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03610_ ), .B1(_03615_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04184_ ) );
AND3_X1 _11466_ ( .A1(_03753_ ), .A2(_00978_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04185_ ) );
AOI21_X1 _11467_ ( .A(_04185_ ), .B1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03532_ ), .ZN(_04186_ ) );
AOI21_X1 _11468_ ( .A(_01049_ ), .B1(_04184_ ), .B2(_04186_ ), .ZN(_04187_ ) );
AOI22_X1 _11469_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03610_ ), .B1(_03615_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04188_ ) );
AND3_X1 _11470_ ( .A1(_03753_ ), .A2(_00978_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04189_ ) );
AOI21_X1 _11471_ ( .A(_04189_ ), .B1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03532_ ), .ZN(_04190_ ) );
AOI21_X1 _11472_ ( .A(_03517_ ), .B1(_04188_ ), .B2(_04190_ ), .ZN(_04191_ ) );
OAI21_X1 _11473_ ( .A(_03641_ ), .B1(_04187_ ), .B2(_04191_ ), .ZN(_04192_ ) );
AND3_X1 _11474_ ( .A1(_00989_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04193_ ) );
AND3_X1 _11475_ ( .A1(_00928_ ), .A2(_00749_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04194_ ) );
OR2_X1 _11476_ ( .A1(_04193_ ), .A2(_04194_ ), .ZN(_04195_ ) );
OAI211_X1 _11477_ ( .A(\u_idu.imm_auipc_lui [20] ), .B(\u_reg.rf[1][2] ), .C1(_02563_ ), .C2(_01078_ ), .ZN(_04196_ ) );
AOI211_X1 _11478_ ( .A(_01049_ ), .B(_04195_ ), .C1(_00956_ ), .C2(_04196_ ), .ZN(_04197_ ) );
OR2_X1 _11479_ ( .A1(_04197_ ), .A2(_00926_ ), .ZN(_04198_ ) );
AOI22_X1 _11480_ ( .A1(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03643_ ), .B1(_03721_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04199_ ) );
AOI21_X1 _11481_ ( .A(_03517_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04200_ ) );
NAND3_X1 _11482_ ( .A1(_03590_ ), .A2(_03560_ ), .A3(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04201_ ) );
AND3_X1 _11483_ ( .A1(_04199_ ), .A2(_04200_ ), .A3(_04201_ ), .ZN(_04202_ ) );
OAI21_X1 _11484_ ( .A(_04192_ ), .B1(_04198_ ), .B2(_04202_ ), .ZN(_04203_ ) );
AOI21_X2 _11485_ ( .A(_03515_ ), .B1(_03508_ ), .B2(_04203_ ), .ZN(_04204_ ) );
OAI21_X1 _11486_ ( .A(_04204_ ), .B1(\ar_data [2] ), .B2(_03509_ ), .ZN(_04205_ ) );
MUX2_X1 _11487_ ( .A(_02675_ ), .B(_04205_ ), .S(_03499_ ), .Z(_04206_ ) );
NOR2_X1 _11488_ ( .A1(_04206_ ), .A2(_03585_ ), .ZN(_04207_ ) );
AOI21_X1 _11489_ ( .A(_04207_ ), .B1(_02362_ ), .B2(_02683_ ), .ZN(_04208_ ) );
AND2_X2 _11490_ ( .A1(_03489_ ), .A2(_03491_ ), .ZN(_04209_ ) );
INV_X2 _11491_ ( .A(_04209_ ), .ZN(_04210_ ) );
OAI21_X2 _11492_ ( .A(_01477_ ), .B1(_04210_ ), .B2(_02683_ ), .ZN(_04211_ ) );
OAI21_X1 _11493_ ( .A(_00744_ ), .B1(_02680_ ), .B2(_02681_ ), .ZN(_04212_ ) );
AND3_X1 _11494_ ( .A1(_01057_ ), .A2(_00745_ ), .A3(_04212_ ), .ZN(_04213_ ) );
AOI221_X1 _11495_ ( .A(_02454_ ), .B1(_01055_ ), .B2(_04208_ ), .C1(_04211_ ), .C2(_04213_ ), .ZN(_00183_ ) );
AND3_X1 _11496_ ( .A1(_02714_ ), .A2(_03974_ ), .A3(_02715_ ), .ZN(_04214_ ) );
NOR2_X1 _11497_ ( .A1(\ar_data [28] ), .A2(_03510_ ), .ZN(_04215_ ) );
AOI22_X1 _11498_ ( .A1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03644_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04216_ ) );
NAND3_X1 _11499_ ( .A1(_03729_ ), .A2(_03543_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04217_ ) );
NAND3_X1 _11500_ ( .A1(_03729_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04218_ ) );
AND4_X1 _11501_ ( .A1(_03519_ ), .A2(_04216_ ), .A3(_04217_ ), .A4(_04218_ ), .ZN(_04219_ ) );
NAND3_X1 _11502_ ( .A1(_03654_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04220_ ) );
NAND3_X1 _11503_ ( .A1(_03605_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04221_ ) );
NAND3_X1 _11504_ ( .A1(_03605_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04222_ ) );
NAND3_X1 _11505_ ( .A1(_04220_ ), .A2(_04221_ ), .A3(_04222_ ), .ZN(_04223_ ) );
AOI211_X1 _11506_ ( .A(_03676_ ), .B(_04223_ ), .C1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03621_ ), .ZN(_04224_ ) );
NOR3_X1 _11507_ ( .A1(_04219_ ), .A2(_04224_ ), .A3(_03660_ ), .ZN(_04225_ ) );
AND3_X1 _11508_ ( .A1(_03606_ ), .A2(_02775_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04226_ ) );
AOI21_X1 _11509_ ( .A(_04226_ ), .B1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03690_ ), .ZN(_04227_ ) );
NAND3_X1 _11510_ ( .A1(_03692_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04228_ ) );
NAND3_X1 _11511_ ( .A1(_03607_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04229_ ) );
NAND4_X1 _11512_ ( .A1(_04227_ ), .A2(_03601_ ), .A3(_04228_ ), .A4(_04229_ ), .ZN(_04230_ ) );
AND2_X1 _11513_ ( .A1(_03528_ ), .A2(\u_reg.rf[1][28] ), .ZN(_04231_ ) );
OAI21_X1 _11514_ ( .A(_03518_ ), .B1(_04231_ ), .B2(_03521_ ), .ZN(_04232_ ) );
AOI221_X4 _11515_ ( .A(_04232_ ), .B1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03612_ ), .C1(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_03722_ ), .ZN(_04233_ ) );
NOR2_X1 _11516_ ( .A1(_04233_ ), .A2(_03641_ ), .ZN(_04234_ ) );
AOI21_X1 _11517_ ( .A(_04225_ ), .B1(_04230_ ), .B2(_04234_ ), .ZN(_04235_ ) );
OAI21_X1 _11518_ ( .A(_03516_ ), .B1(_03507_ ), .B2(_04235_ ), .ZN(_04236_ ) );
OR2_X2 _11519_ ( .A1(_04215_ ), .A2(_04236_ ), .ZN(_04237_ ) );
AOI211_X1 _11520_ ( .A(_03586_ ), .B(_04214_ ), .C1(_04237_ ), .C2(_03629_ ), .ZN(_04238_ ) );
AND2_X1 _11521_ ( .A1(_02722_ ), .A2(_02568_ ), .ZN(_04239_ ) );
OAI21_X1 _11522_ ( .A(_03998_ ), .B1(_04238_ ), .B2(_04239_ ), .ZN(_04240_ ) );
NAND2_X1 _11523_ ( .A1(_03498_ ), .A2(_04240_ ), .ZN(_00184_ ) );
OAI211_X1 _11524_ ( .A(_01070_ ), .B(_02779_ ), .C1(_03945_ ), .C2(_03946_ ), .ZN(_04241_ ) );
NAND4_X1 _11525_ ( .A1(_02509_ ), .A2(_02765_ ), .A3(_01597_ ), .A4(_01381_ ), .ZN(_04242_ ) );
AND3_X1 _11526_ ( .A1(_02763_ ), .A2(_03974_ ), .A3(_04242_ ), .ZN(_04243_ ) );
AOI21_X1 _11527_ ( .A(_03623_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04244_ ) );
NAND3_X1 _11528_ ( .A1(_03607_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04245_ ) );
NAND3_X1 _11529_ ( .A1(_04095_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04246_ ) );
NAND3_X1 _11530_ ( .A1(_03680_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04247_ ) );
NAND4_X1 _11531_ ( .A1(_04244_ ), .A2(_04245_ ), .A3(_04246_ ), .A4(_04247_ ), .ZN(_04248_ ) );
AOI21_X1 _11532_ ( .A(_03677_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04249_ ) );
NAND3_X1 _11533_ ( .A1(_03680_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04250_ ) );
NAND3_X1 _11534_ ( .A1(_04095_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04251_ ) );
NAND3_X1 _11535_ ( .A1(_03680_ ), .A2(fanout_net_21 ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04252_ ) );
NAND4_X1 _11536_ ( .A1(_04249_ ), .A2(_04250_ ), .A3(_04251_ ), .A4(_04252_ ), .ZN(_04253_ ) );
NAND3_X1 _11537_ ( .A1(_04248_ ), .A2(_04253_ ), .A3(_03687_ ), .ZN(_04254_ ) );
AND3_X1 _11538_ ( .A1(_03549_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04255_ ) );
AOI221_X4 _11539_ ( .A(_04255_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03553_ ), .ZN(_04256_ ) );
NAND3_X1 _11540_ ( .A1(_03692_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04257_ ) );
AND3_X1 _11541_ ( .A1(_04256_ ), .A2(_03557_ ), .A3(_04257_ ), .ZN(_04258_ ) );
AND3_X1 _11542_ ( .A1(_03541_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04259_ ) );
AOI21_X1 _11543_ ( .A(_04259_ ), .B1(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03672_ ), .ZN(_04260_ ) );
AOI211_X1 _11544_ ( .A(_03562_ ), .B(_02748_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_04261_ ) );
OAI211_X1 _11545_ ( .A(_04260_ ), .B(_03678_ ), .C1(_03559_ ), .C2(_04261_ ), .ZN(_04262_ ) );
NAND2_X1 _11546_ ( .A1(_04262_ ), .A2(_03661_ ), .ZN(_04263_ ) );
OAI21_X1 _11547_ ( .A(_04254_ ), .B1(_04258_ ), .B2(_04263_ ), .ZN(_04264_ ) );
AOI21_X2 _11548_ ( .A(_03669_ ), .B1(_03511_ ), .B2(_04264_ ), .ZN(_04265_ ) );
OAI21_X1 _11549_ ( .A(_04265_ ), .B1(\ar_data [1] ), .B2(_03704_ ), .ZN(_04266_ ) );
AOI211_X1 _11550_ ( .A(_03973_ ), .B(_04243_ ), .C1(_04266_ ), .C2(_03994_ ), .ZN(_04267_ ) );
NOR2_X1 _11551_ ( .A1(_02778_ ), .A2(_03631_ ), .ZN(_04268_ ) );
OAI21_X1 _11552_ ( .A(_03998_ ), .B1(_04267_ ), .B2(_04268_ ), .ZN(_04269_ ) );
NAND2_X1 _11553_ ( .A1(_04241_ ), .A2(_04269_ ), .ZN(_00185_ ) );
AOI22_X1 _11554_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03637_ ), .B1(_03615_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04270_ ) );
AOI22_X1 _11555_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03552_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04271_ ) );
AOI21_X1 _11556_ ( .A(_03555_ ), .B1(_04270_ ), .B2(_04271_ ), .ZN(_04272_ ) );
AND3_X1 _11557_ ( .A1(_03527_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04273_ ) );
AOI21_X1 _11558_ ( .A(_04273_ ), .B1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03611_ ), .ZN(_04274_ ) );
AOI22_X1 _11559_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03643_ ), .B1(_03619_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04275_ ) );
AOI21_X1 _11560_ ( .A(_03675_ ), .B1(_04274_ ), .B2(_04275_ ), .ZN(_04276_ ) );
OAI21_X1 _11561_ ( .A(_03641_ ), .B1(_04272_ ), .B2(_04276_ ), .ZN(_04277_ ) );
AND3_X1 _11562_ ( .A1(_03520_ ), .A2(_03560_ ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04278_ ) );
AOI21_X1 _11563_ ( .A(_04278_ ), .B1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03721_ ), .ZN(_04279_ ) );
AOI211_X1 _11564_ ( .A(_03560_ ), .B(_02787_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_04280_ ) );
OAI211_X1 _11565_ ( .A(_04279_ ), .B(_03518_ ), .C1(_03654_ ), .C2(_04280_ ), .ZN(_04281_ ) );
AOI22_X1 _11566_ ( .A1(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03552_ ), .B1(_03721_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04282_ ) );
AOI21_X1 _11567_ ( .A(_03675_ ), .B1(_03533_ ), .B2(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04283_ ) );
NAND3_X1 _11568_ ( .A1(_03590_ ), .A2(_03523_ ), .A3(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04284_ ) );
NAND3_X1 _11569_ ( .A1(_04282_ ), .A2(_04283_ ), .A3(_04284_ ), .ZN(_04285_ ) );
NAND3_X1 _11570_ ( .A1(_04281_ ), .A2(_03537_ ), .A3(_04285_ ), .ZN(_04286_ ) );
AND2_X1 _11571_ ( .A1(_04277_ ), .A2(_04286_ ), .ZN(_04287_ ) );
OR2_X1 _11572_ ( .A1(_03507_ ), .A2(_04287_ ), .ZN(_04288_ ) );
AND2_X1 _11573_ ( .A1(_02809_ ), .A2(_02811_ ), .ZN(\ar_data [0] ) );
OAI211_X1 _11574_ ( .A(_04288_ ), .B(_03516_ ), .C1(\ar_data [0] ), .C2(_03710_ ), .ZN(_04289_ ) );
AOI21_X1 _11575_ ( .A(_03585_ ), .B1(_04289_ ), .B2(_03499_ ), .ZN(_04290_ ) );
NAND4_X1 _11576_ ( .A1(_02509_ ), .A2(_02820_ ), .A3(_01444_ ), .A4(_01381_ ), .ZN(_04291_ ) );
OAI211_X1 _11577_ ( .A(_03579_ ), .B(_04291_ ), .C1(_02818_ ), .C2(_02492_ ), .ZN(_04292_ ) );
AOI22_X1 _11578_ ( .A1(_04290_ ), .A2(_04292_ ), .B1(_01490_ ), .B2(_02830_ ), .ZN(_04293_ ) );
NAND4_X1 _11579_ ( .A1(_03489_ ), .A2(_01475_ ), .A3(_02830_ ), .A4(_03491_ ), .ZN(_04294_ ) );
AND3_X1 _11580_ ( .A1(_00717_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(_00718_ ), .ZN(_04295_ ) );
AOI21_X1 _11581_ ( .A(_04295_ ), .B1(_03739_ ), .B2(_03740_ ), .ZN(_04296_ ) );
AOI221_X1 _11582_ ( .A(_02454_ ), .B1(_01055_ ), .B2(_04293_ ), .C1(_04294_ ), .C2(_04296_ ), .ZN(_00186_ ) );
AND3_X1 _11583_ ( .A1(_02859_ ), .A2(_03974_ ), .A3(_02860_ ), .ZN(_04297_ ) );
AOI22_X1 _11584_ ( .A1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03553_ ), .B1(_03534_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04298_ ) );
NAND3_X1 _11585_ ( .A1(_03655_ ), .A2(_03562_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04299_ ) );
NAND3_X1 _11586_ ( .A1(_03655_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04300_ ) );
AND4_X1 _11587_ ( .A1(_03519_ ), .A2(_04298_ ), .A3(_04299_ ), .A4(_04300_ ), .ZN(_04301_ ) );
NAND3_X1 _11588_ ( .A1(_03522_ ), .A2(_03543_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04302_ ) );
NAND3_X1 _11589_ ( .A1(_03529_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04303_ ) );
NAND3_X1 _11590_ ( .A1(_03529_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04304_ ) );
NAND3_X1 _11591_ ( .A1(_04302_ ), .A2(_04303_ ), .A3(_04304_ ), .ZN(_04305_ ) );
AOI211_X1 _11592_ ( .A(_03519_ ), .B(_04305_ ), .C1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03535_ ), .ZN(_04306_ ) );
OR3_X1 _11593_ ( .A1(_04301_ ), .A2(_04306_ ), .A3(_03538_ ), .ZN(_04307_ ) );
AND3_X1 _11594_ ( .A1(_03549_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04308_ ) );
AOI221_X4 _11595_ ( .A(_04308_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03553_ ), .ZN(_04309_ ) );
NAND3_X1 _11596_ ( .A1(_03559_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04310_ ) );
NAND3_X1 _11597_ ( .A1(_04309_ ), .A2(_03557_ ), .A3(_04310_ ), .ZN(_04311_ ) );
AND3_X1 _11598_ ( .A1(_03541_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04312_ ) );
AOI21_X1 _11599_ ( .A(_04312_ ), .B1(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03672_ ), .ZN(_04313_ ) );
AND2_X1 _11600_ ( .A1(_03571_ ), .A2(\u_reg.rf[1][27] ), .ZN(_04314_ ) );
OAI211_X1 _11601_ ( .A(_04313_ ), .B(_03678_ ), .C1(_03559_ ), .C2(_04314_ ), .ZN(_04315_ ) );
NAND3_X1 _11602_ ( .A1(_04311_ ), .A2(_03661_ ), .A3(_04315_ ), .ZN(_04316_ ) );
NAND2_X1 _11603_ ( .A1(_04307_ ), .A2(_04316_ ), .ZN(_04317_ ) );
AOI21_X1 _11604_ ( .A(_03670_ ), .B1(_03671_ ), .B2(_04317_ ), .ZN(_04318_ ) );
OAI21_X1 _11605_ ( .A(_04318_ ), .B1(\ar_data [27] ), .B2(_03704_ ), .ZN(_04319_ ) );
AOI211_X1 _11606_ ( .A(_03973_ ), .B(_04297_ ), .C1(_04319_ ), .C2(_03994_ ), .ZN(_04320_ ) );
NOR2_X1 _11607_ ( .A1(_02865_ ), .A2(_03631_ ), .ZN(_04321_ ) );
OAI21_X1 _11608_ ( .A(_03998_ ), .B1(_04320_ ), .B2(_04321_ ), .ZN(_04322_ ) );
NAND2_X1 _11609_ ( .A1(_03498_ ), .A2(_04322_ ), .ZN(_00187_ ) );
NAND2_X1 _11610_ ( .A1(_01596_ ), .A2(_01597_ ), .ZN(_04323_ ) );
AOI21_X1 _11611_ ( .A(_04323_ ), .B1(_00841_ ), .B2(_00842_ ), .ZN(_04324_ ) );
NOR3_X1 _11612_ ( .A1(_02896_ ), .A2(_03500_ ), .A3(_04324_ ), .ZN(_04325_ ) );
NOR2_X2 _11613_ ( .A1(\ar_data [26] ), .A2(_03510_ ), .ZN(_04326_ ) );
AOI22_X1 _11614_ ( .A1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03553_ ), .B1(_03612_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04327_ ) );
AOI21_X1 _11615_ ( .A(_03539_ ), .B1(_03534_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04328_ ) );
NAND3_X1 _11616_ ( .A1(_03606_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04329_ ) );
AND3_X1 _11617_ ( .A1(_04327_ ), .A2(_04328_ ), .A3(_04329_ ), .ZN(_04330_ ) );
NAND3_X1 _11618_ ( .A1(_03605_ ), .A2(_02774_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04331_ ) );
NAND2_X1 _11619_ ( .A1(_04331_ ), .A2(_03539_ ), .ZN(_04332_ ) );
NAND3_X1 _11620_ ( .A1(_03654_ ), .A2(_03524_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04333_ ) );
NAND3_X1 _11621_ ( .A1(_03605_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04334_ ) );
NAND2_X1 _11622_ ( .A1(_04333_ ), .A2(_04334_ ), .ZN(_04335_ ) );
AOI211_X1 _11623_ ( .A(_04332_ ), .B(_04335_ ), .C1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03621_ ), .ZN(_04336_ ) );
NOR3_X1 _11624_ ( .A1(_04330_ ), .A2(_04336_ ), .A3(_03660_ ), .ZN(_04337_ ) );
AOI21_X1 _11625_ ( .A(_03677_ ), .B1(_03690_ ), .B2(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04338_ ) );
NAND3_X1 _11626_ ( .A1(_03692_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04339_ ) );
NAND3_X1 _11627_ ( .A1(_03607_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04340_ ) );
NAND3_X1 _11628_ ( .A1(_03607_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04341_ ) );
NAND4_X1 _11629_ ( .A1(_04338_ ), .A2(_04339_ ), .A3(_04340_ ), .A4(_04341_ ), .ZN(_04342_ ) );
AND3_X1 _11630_ ( .A1(_03549_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04343_ ) );
AOI21_X1 _11631_ ( .A(_04343_ ), .B1(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B2(_03613_ ), .ZN(_04344_ ) );
AND2_X1 _11632_ ( .A1(_03541_ ), .A2(\u_reg.rf[1][26] ), .ZN(_04345_ ) );
OAI211_X1 _11633_ ( .A(_04344_ ), .B(_03677_ ), .C1(_04095_ ), .C2(_04345_ ), .ZN(_04346_ ) );
AND2_X1 _11634_ ( .A1(_04346_ ), .A2(_03538_ ), .ZN(_04347_ ) );
AOI21_X1 _11635_ ( .A(_04337_ ), .B1(_04342_ ), .B2(_04347_ ), .ZN(_04348_ ) );
OAI21_X1 _11636_ ( .A(_03516_ ), .B1(_03507_ ), .B2(_04348_ ), .ZN(_04349_ ) );
OR2_X2 _11637_ ( .A1(_04326_ ), .A2(_04349_ ), .ZN(_04350_ ) );
AOI211_X1 _11638_ ( .A(_03973_ ), .B(_04325_ ), .C1(_04350_ ), .C2(_03994_ ), .ZN(_04351_ ) );
NOR2_X1 _11639_ ( .A1(_02904_ ), .A2(_03631_ ), .ZN(_04352_ ) );
OAI21_X1 _11640_ ( .A(_03998_ ), .B1(_04351_ ), .B2(_04352_ ), .ZN(_04353_ ) );
NAND2_X1 _11641_ ( .A1(_03498_ ), .A2(_04353_ ), .ZN(_00188_ ) );
AND3_X1 _11642_ ( .A1(_02933_ ), .A2(_03974_ ), .A3(_02934_ ), .ZN(_04354_ ) );
AOI22_X1 _11643_ ( .A1(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04355_ ) );
NAND3_X1 _11644_ ( .A1(_03692_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04356_ ) );
NAND3_X1 _11645_ ( .A1(_03692_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04357_ ) );
NAND4_X1 _11646_ ( .A1(_04355_ ), .A2(_03678_ ), .A3(_04356_ ), .A4(_04357_ ), .ZN(_04358_ ) );
AOI21_X1 _11647_ ( .A(_03677_ ), .B1(_03673_ ), .B2(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04359_ ) );
NAND3_X1 _11648_ ( .A1(_03692_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04360_ ) );
NAND3_X1 _11649_ ( .A1(_03680_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04361_ ) );
NAND3_X1 _11650_ ( .A1(_03680_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04362_ ) );
NAND4_X1 _11651_ ( .A1(_04359_ ), .A2(_04360_ ), .A3(_04361_ ), .A4(_04362_ ), .ZN(_04363_ ) );
NAND3_X1 _11652_ ( .A1(_04358_ ), .A2(_03687_ ), .A3(_04363_ ), .ZN(_04364_ ) );
AND3_X1 _11653_ ( .A1(_03655_ ), .A2(_03562_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04365_ ) );
AND3_X1 _11654_ ( .A1(_03729_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04366_ ) );
AOI21_X1 _11655_ ( .A(_03655_ ), .B1(\u_reg.rf[1][25] ), .B2(_03606_ ), .ZN(_04367_ ) );
NOR3_X1 _11656_ ( .A1(_04365_ ), .A2(_04366_ ), .A3(_04367_ ), .ZN(_04368_ ) );
NAND3_X1 _11657_ ( .A1(_03729_ ), .A2(_03543_ ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04369_ ) );
NAND3_X1 _11658_ ( .A1(_03729_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04370_ ) );
NAND2_X1 _11659_ ( .A1(_04369_ ), .A2(_04370_ ), .ZN(_04371_ ) );
MUX2_X1 _11660_ ( .A(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03529_ ), .Z(_04372_ ) );
AOI21_X1 _11661_ ( .A(_04371_ ), .B1(_04372_ ), .B2(_03567_ ), .ZN(_04373_ ) );
MUX2_X1 _11662_ ( .A(_04368_ ), .B(_04373_ ), .S(_03601_ ), .Z(_04374_ ) );
OAI21_X1 _11663_ ( .A(_04364_ ), .B1(_04374_ ), .B2(_03687_ ), .ZN(_04375_ ) );
AOI21_X1 _11664_ ( .A(_03670_ ), .B1(_03671_ ), .B2(_04375_ ), .ZN(_04376_ ) );
OAI21_X2 _11665_ ( .A(_04376_ ), .B1(\ar_data [25] ), .B2(_03704_ ), .ZN(_04377_ ) );
AOI211_X1 _11666_ ( .A(_03973_ ), .B(_04354_ ), .C1(_04377_ ), .C2(_03994_ ), .ZN(_04378_ ) );
AND2_X1 _11667_ ( .A1(_02939_ ), .A2(_02568_ ), .ZN(_04379_ ) );
OAI21_X1 _11668_ ( .A(_03998_ ), .B1(_04378_ ), .B2(_04379_ ), .ZN(_04380_ ) );
NAND2_X1 _11669_ ( .A1(_03498_ ), .A2(_04380_ ), .ZN(_00189_ ) );
NAND3_X1 _11670_ ( .A1(_02977_ ), .A2(_03580_ ), .A3(_02978_ ), .ZN(_04381_ ) );
OR2_X2 _11671_ ( .A1(\ar_data [24] ), .A2(_03710_ ), .ZN(_04382_ ) );
AND3_X1 _11672_ ( .A1(_03521_ ), .A2(_03561_ ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04383_ ) );
AOI21_X1 _11673_ ( .A(_04383_ ), .B1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03929_ ), .ZN(_04384_ ) );
AOI22_X1 _11674_ ( .A1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03553_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04385_ ) );
AND3_X1 _11675_ ( .A1(_04384_ ), .A2(_04385_ ), .A3(_03556_ ), .ZN(_04386_ ) );
AOI21_X1 _11676_ ( .A(_03601_ ), .B1(_03690_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04387_ ) );
AND3_X1 _11677_ ( .A1(_03549_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04388_ ) );
AOI221_X4 _11678_ ( .A(_04388_ ), .B1(_03644_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03613_ ), .ZN(_04389_ ) );
AOI211_X1 _11679_ ( .A(_03661_ ), .B(_04386_ ), .C1(_04387_ ), .C2(_04389_ ), .ZN(_04390_ ) );
AOI22_X1 _11680_ ( .A1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03553_ ), .B1(_03929_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04391_ ) );
AOI21_X1 _11681_ ( .A(_03676_ ), .B1(_03621_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04392_ ) );
NAND3_X1 _11682_ ( .A1(_03558_ ), .A2(_03569_ ), .A3(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04393_ ) );
NAND3_X1 _11683_ ( .A1(_04391_ ), .A2(_04392_ ), .A3(_04393_ ), .ZN(_04394_ ) );
AOI22_X1 _11684_ ( .A1(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_03613_ ), .B1(_03929_ ), .B2(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04395_ ) );
OAI21_X1 _11685_ ( .A(_03567_ ), .B1(_00958_ ), .B2(_02958_ ), .ZN(_04396_ ) );
NAND3_X1 _11686_ ( .A1(_04395_ ), .A2(_03677_ ), .A3(_04396_ ), .ZN(_04397_ ) );
AND3_X1 _11687_ ( .A1(_04394_ ), .A2(_04397_ ), .A3(_03538_ ), .ZN(_04398_ ) );
OAI21_X1 _11688_ ( .A(_03510_ ), .B1(_04390_ ), .B2(_04398_ ), .ZN(_04399_ ) );
AND3_X2 _11689_ ( .A1(_04382_ ), .A2(_03516_ ), .A3(_04399_ ), .ZN(_04400_ ) );
OAI211_X1 _11690_ ( .A(_03578_ ), .B(_04381_ ), .C1(_04400_ ), .C2(_03580_ ), .ZN(_04401_ ) );
OAI21_X1 _11691_ ( .A(_04401_ ), .B1(_03631_ ), .B2(_02983_ ), .ZN(_04402_ ) );
NAND2_X1 _11692_ ( .A1(_04402_ ), .A2(_00302_ ), .ZN(_04403_ ) );
NAND2_X1 _11693_ ( .A1(_03498_ ), .A2(_04403_ ), .ZN(_00190_ ) );
AOI21_X1 _11694_ ( .A(_04323_ ), .B1(_00847_ ), .B2(_00848_ ), .ZN(_04404_ ) );
NOR3_X1 _11695_ ( .A1(_03022_ ), .A2(_03500_ ), .A3(_04404_ ), .ZN(_04405_ ) );
AND3_X1 _11696_ ( .A1(_03520_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04406_ ) );
AOI221_X4 _11697_ ( .A(_04406_ ), .B1(_03643_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03611_ ), .ZN(_04407_ ) );
AOI21_X1 _11698_ ( .A(_03555_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04408_ ) );
AOI21_X1 _11699_ ( .A(_03676_ ), .B1(_03534_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04409_ ) );
AND3_X1 _11700_ ( .A1(_03527_ ), .A2(_02773_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04410_ ) );
AOI221_X4 _11701_ ( .A(_04410_ ), .B1(_03721_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_03637_ ), .ZN(_04411_ ) );
AOI221_X4 _11702_ ( .A(_03660_ ), .B1(_04407_ ), .B2(_04408_ ), .C1(_04409_ ), .C2(_04411_ ), .ZN(_04412_ ) );
AND3_X1 _11703_ ( .A1(_03548_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04413_ ) );
AOI221_X4 _11704_ ( .A(_04413_ ), .B1(_03533_ ), .B2(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03552_ ), .ZN(_04414_ ) );
NAND3_X1 _11705_ ( .A1(_03655_ ), .A2(_03562_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04415_ ) );
NAND3_X1 _11706_ ( .A1(_04414_ ), .A2(_03623_ ), .A3(_04415_ ), .ZN(_04416_ ) );
AND3_X1 _11707_ ( .A1(_03521_ ), .A2(_03561_ ), .A3(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04417_ ) );
AOI21_X1 _11708_ ( .A(_04417_ ), .B1(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03929_ ), .ZN(_04418_ ) );
AOI211_X1 _11709_ ( .A(_03524_ ), .B(_03003_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_04419_ ) );
OAI211_X1 _11710_ ( .A(_04418_ ), .B(_03519_ ), .C1(_04095_ ), .C2(_04419_ ), .ZN(_04420_ ) );
AND3_X1 _11711_ ( .A1(_04416_ ), .A2(_03538_ ), .A3(_04420_ ), .ZN(_04421_ ) );
OR2_X1 _11712_ ( .A1(_04412_ ), .A2(_04421_ ), .ZN(_04422_ ) );
AOI21_X1 _11713_ ( .A(_03670_ ), .B1(_03511_ ), .B2(_04422_ ), .ZN(_04423_ ) );
OAI21_X2 _11714_ ( .A(_04423_ ), .B1(\ar_data [23] ), .B2(_03704_ ), .ZN(_04424_ ) );
AOI211_X1 _11715_ ( .A(_03973_ ), .B(_04405_ ), .C1(_04424_ ), .C2(_03994_ ), .ZN(_04425_ ) );
NOR2_X1 _11716_ ( .A1(_03030_ ), .A2(_03631_ ), .ZN(_04426_ ) );
OAI21_X1 _11717_ ( .A(_03998_ ), .B1(_04425_ ), .B2(_04426_ ), .ZN(_04427_ ) );
NAND2_X1 _11718_ ( .A1(_03497_ ), .A2(_04427_ ), .ZN(_00191_ ) );
AND3_X1 _11719_ ( .A1(_03069_ ), .A2(_03974_ ), .A3(_03070_ ), .ZN(_04428_ ) );
AOI22_X1 _11720_ ( .A1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_03684_ ), .B1(_03535_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04429_ ) );
NAND3_X1 _11721_ ( .A1(_04095_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04430_ ) );
NAND3_X1 _11722_ ( .A1(_04095_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04431_ ) );
NAND4_X1 _11723_ ( .A1(_04429_ ), .A2(_03677_ ), .A3(_04430_ ), .A4(_04431_ ), .ZN(_04432_ ) );
OAI21_X1 _11724_ ( .A(_03601_ ), .B1(_04085_ ), .B2(_03046_ ), .ZN(_04433_ ) );
NAND3_X1 _11725_ ( .A1(_03692_ ), .A2(_04096_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04434_ ) );
NAND3_X1 _11726_ ( .A1(_04095_ ), .A2(\u_idu.imm_auipc_lui [20] ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04435_ ) );
NAND3_X1 _11727_ ( .A1(_03680_ ), .A2(_02776_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04436_ ) );
NAND3_X1 _11728_ ( .A1(_04434_ ), .A2(_04435_ ), .A3(_04436_ ), .ZN(_04437_ ) );
OAI211_X1 _11729_ ( .A(_04432_ ), .B(_03687_ ), .C1(_04433_ ), .C2(_04437_ ), .ZN(_04438_ ) );
AND3_X1 _11730_ ( .A1(_03549_ ), .A2(\u_idu.imm_auipc_lui [21] ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04439_ ) );
AOI221_X4 _11731_ ( .A(_04439_ ), .B1(_03551_ ), .B2(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_03553_ ), .ZN(_04440_ ) );
NAND3_X1 _11732_ ( .A1(_03559_ ), .A2(_03563_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04441_ ) );
NAND3_X1 _11733_ ( .A1(_04440_ ), .A2(_03557_ ), .A3(_04441_ ), .ZN(_04442_ ) );
AND3_X1 _11734_ ( .A1(_03729_ ), .A2(_03543_ ), .A3(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04443_ ) );
AOI21_X1 _11735_ ( .A(_04443_ ), .B1(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_03929_ ), .ZN(_04444_ ) );
AOI211_X1 _11736_ ( .A(_03569_ ), .B(_03058_ ), .C1(_00921_ ), .C2(_00923_ ), .ZN(_04445_ ) );
OAI211_X1 _11737_ ( .A(_04444_ ), .B(_03678_ ), .C1(_03559_ ), .C2(_04445_ ), .ZN(_04446_ ) );
NAND2_X1 _11738_ ( .A1(_04442_ ), .A2(_04446_ ), .ZN(_04447_ ) );
OAI21_X1 _11739_ ( .A(_04438_ ), .B1(_04447_ ), .B2(_03687_ ), .ZN(_04448_ ) );
AOI21_X1 _11740_ ( .A(_03670_ ), .B1(_03511_ ), .B2(_04448_ ), .ZN(_04449_ ) );
OAI21_X1 _11741_ ( .A(_04449_ ), .B1(\ar_data [22] ), .B2(_03704_ ), .ZN(_04450_ ) );
AOI211_X1 _11742_ ( .A(_03973_ ), .B(_04428_ ), .C1(_04450_ ), .C2(_03994_ ), .ZN(_04451_ ) );
NOR2_X1 _11743_ ( .A1(_03075_ ), .A2(_03631_ ), .ZN(_04452_ ) );
OAI21_X1 _11744_ ( .A(_01569_ ), .B1(_04451_ ), .B2(_04452_ ), .ZN(_04453_ ) );
NAND2_X1 _11745_ ( .A1(_03497_ ), .A2(_04453_ ), .ZN(_00192_ ) );
BUF_X2 _11746_ ( .A(_00862_ ), .Z(_04454_ ) );
AND3_X1 _11747_ ( .A1(_00920_ ), .A2(_00866_ ), .A3(_04454_ ), .ZN(_00193_ ) );
BUF_X4 _11748_ ( .A(_00880_ ), .Z(_04455_ ) );
BUF_X4 _11749_ ( .A(_00855_ ), .Z(_04456_ ) );
NOR3_X1 _11750_ ( .A1(_00905_ ), .A2(_04455_ ), .A3(_04456_ ), .ZN(_00194_ ) );
NOR3_X1 _11751_ ( .A1(_00910_ ), .A2(_04455_ ), .A3(_04456_ ), .ZN(_00195_ ) );
NOR3_X1 _11752_ ( .A1(_00914_ ), .A2(_04455_ ), .A3(_00882_ ), .ZN(_00196_ ) );
AOI21_X1 _11753_ ( .A(_02456_ ), .B1(_01470_ ), .B2(_01473_ ), .ZN(_00197_ ) );
AOI21_X1 _11754_ ( .A(_02456_ ), .B1(_01595_ ), .B2(_01598_ ), .ZN(_00198_ ) );
AOI21_X1 _11755_ ( .A(_02456_ ), .B1(_01658_ ), .B2(_01659_ ), .ZN(_00199_ ) );
AOI21_X1 _11756_ ( .A(_02456_ ), .B1(_01714_ ), .B2(_01716_ ), .ZN(_00200_ ) );
AOI21_X1 _11757_ ( .A(_02456_ ), .B1(_01773_ ), .B2(_01775_ ), .ZN(_00201_ ) );
AOI21_X1 _11758_ ( .A(_02456_ ), .B1(_01840_ ), .B2(_01841_ ), .ZN(_00202_ ) );
AOI21_X1 _11759_ ( .A(_02456_ ), .B1(_01896_ ), .B2(_01897_ ), .ZN(_00203_ ) );
AOI21_X1 _11760_ ( .A(_02456_ ), .B1(_01948_ ), .B2(_01949_ ), .ZN(_00204_ ) );
AOI21_X1 _11761_ ( .A(_02456_ ), .B1(_01986_ ), .B2(_01987_ ), .ZN(_00205_ ) );
BUF_X4 _11762_ ( .A(_02455_ ), .Z(_04457_ ) );
AOI21_X1 _11763_ ( .A(_04457_ ), .B1(_02042_ ), .B2(_02043_ ), .ZN(_00206_ ) );
AOI21_X1 _11764_ ( .A(_04457_ ), .B1(_02089_ ), .B2(_02090_ ), .ZN(_00207_ ) );
AOI21_X1 _11765_ ( .A(_04457_ ), .B1(_02131_ ), .B2(_02136_ ), .ZN(_00208_ ) );
AOI21_X1 _11766_ ( .A(_04457_ ), .B1(_02171_ ), .B2(_02172_ ), .ZN(_00209_ ) );
AOI21_X1 _11767_ ( .A(_04457_ ), .B1(_02211_ ), .B2(_02217_ ), .ZN(_00210_ ) );
AOI21_X1 _11768_ ( .A(_04457_ ), .B1(_02265_ ), .B2(_02266_ ), .ZN(_00211_ ) );
AOI21_X1 _11769_ ( .A(_04457_ ), .B1(_02311_ ), .B2(_02312_ ), .ZN(_00212_ ) );
AOI21_X1 _11770_ ( .A(_04457_ ), .B1(_02352_ ), .B2(_02353_ ), .ZN(_00213_ ) );
AOI21_X1 _11771_ ( .A(_04457_ ), .B1(_02396_ ), .B2(_02397_ ), .ZN(_00214_ ) );
AOI21_X1 _11772_ ( .A(_04457_ ), .B1(_02447_ ), .B2(_02448_ ), .ZN(_00215_ ) );
AND3_X1 _11773_ ( .A1(_01596_ ), .A2(_02500_ ), .A3(_01597_ ), .ZN(_04458_ ) );
NOR2_X1 _11774_ ( .A1(_02499_ ), .A2(_04458_ ), .ZN(_04459_ ) );
BUF_X4 _11775_ ( .A(_02454_ ), .Z(_04460_ ) );
BUF_X4 _11776_ ( .A(_04460_ ), .Z(_04461_ ) );
NOR2_X1 _11777_ ( .A1(_04459_ ), .A2(_04461_ ), .ZN(_00216_ ) );
BUF_X4 _11778_ ( .A(_02455_ ), .Z(_04462_ ) );
AOI21_X1 _11779_ ( .A(_04462_ ), .B1(_02556_ ), .B2(_02557_ ), .ZN(_00217_ ) );
AOI21_X1 _11780_ ( .A(_04462_ ), .B1(_02609_ ), .B2(_02610_ ), .ZN(_00218_ ) );
NOR2_X1 _11781_ ( .A1(_02675_ ), .A2(_04461_ ), .ZN(_00219_ ) );
AOI21_X1 _11782_ ( .A(_04462_ ), .B1(_02714_ ), .B2(_02715_ ), .ZN(_00220_ ) );
AOI21_X1 _11783_ ( .A(_04462_ ), .B1(_02763_ ), .B2(_04242_ ), .ZN(_00221_ ) );
NOR2_X1 _11784_ ( .A1(_02822_ ), .A2(_04461_ ), .ZN(_00222_ ) );
AOI21_X1 _11785_ ( .A(_04462_ ), .B1(_02859_ ), .B2(_02860_ ), .ZN(_00223_ ) );
NOR2_X1 _11786_ ( .A1(_02898_ ), .A2(_04461_ ), .ZN(_00224_ ) );
AOI21_X1 _11787_ ( .A(_04462_ ), .B1(_02933_ ), .B2(_02934_ ), .ZN(_00225_ ) );
AOI21_X1 _11788_ ( .A(_04462_ ), .B1(_02977_ ), .B2(_02978_ ), .ZN(_00226_ ) );
NOR2_X1 _11789_ ( .A1(_03024_ ), .A2(_04461_ ), .ZN(_00227_ ) );
AOI21_X1 _11790_ ( .A(_04462_ ), .B1(_03069_ ), .B2(_03070_ ), .ZN(_00228_ ) );
NOR3_X1 _11791_ ( .A1(_01100_ ), .A2(_04456_ ), .A3(_04455_ ), .ZN(_00232_ ) );
NOR3_X1 _11792_ ( .A1(flush_$_OR__Y_B ), .A2(_01104_ ), .A3(_00882_ ), .ZN(_00233_ ) );
NOR2_X1 _11793_ ( .A1(_00723_ ), .A2(_04461_ ), .ZN(_00234_ ) );
AND3_X1 _11794_ ( .A1(_00864_ ), .A2(\de_pc [31] ), .A3(_00866_ ), .ZN(_00235_ ) );
NOR4_X1 _11795_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_01508_ ), .ZN(_00236_ ) );
AND3_X1 _11796_ ( .A1(_00864_ ), .A2(\de_pc [21] ), .A3(_00866_ ), .ZN(_00237_ ) );
AND3_X1 _11797_ ( .A1(_00864_ ), .A2(\de_pc [20] ), .A3(_00866_ ), .ZN(_00238_ ) );
AND3_X1 _11798_ ( .A1(_00864_ ), .A2(\de_pc [19] ), .A3(_00866_ ), .ZN(_00239_ ) );
NOR4_X1 _11799_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_01844_ ), .ZN(_00240_ ) );
NOR4_X1 _11800_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_01899_ ), .ZN(_00241_ ) );
AND3_X1 _11801_ ( .A1(_00864_ ), .A2(\de_pc [16] ), .A3(_00866_ ), .ZN(_00242_ ) );
NOR4_X1 _11802_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_00885_ ), .A4(_01989_ ), .ZN(_00243_ ) );
BUF_X4 _11803_ ( .A(_00858_ ), .Z(_04463_ ) );
NOR4_X1 _11804_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_04463_ ), .A4(_02045_ ), .ZN(_00244_ ) );
NOR4_X1 _11805_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_04463_ ), .A4(_02092_ ), .ZN(_00245_ ) );
AND3_X1 _11806_ ( .A1(_00864_ ), .A2(\de_pc [12] ), .A3(_00866_ ), .ZN(_00246_ ) );
CLKBUF_X2 _11807_ ( .A(_00865_ ), .Z(_04464_ ) );
AND3_X1 _11808_ ( .A1(_00864_ ), .A2(\de_pc [29] ), .A3(_04464_ ), .ZN(_00247_ ) );
NOR4_X1 _11809_ ( .A1(_00889_ ), .A2(fanout_net_1 ), .A3(_04463_ ), .A4(_02219_ ), .ZN(_00248_ ) );
AND3_X1 _11810_ ( .A1(_00864_ ), .A2(\de_pc [10] ), .A3(_04464_ ), .ZN(_00249_ ) );
AND3_X1 _11811_ ( .A1(_00864_ ), .A2(\de_pc [9] ), .A3(_04464_ ), .ZN(_00250_ ) );
NOR4_X1 _11812_ ( .A1(_00889_ ), .A2(fanout_net_2 ), .A3(_04463_ ), .A4(_02355_ ), .ZN(_00251_ ) );
CLKBUF_X2 _11813_ ( .A(_00863_ ), .Z(_04465_ ) );
AND3_X1 _11814_ ( .A1(_04465_ ), .A2(\de_pc [7] ), .A3(_04464_ ), .ZN(_00252_ ) );
AND3_X1 _11815_ ( .A1(_04465_ ), .A2(\de_pc [6] ), .A3(_04464_ ), .ZN(_00253_ ) );
NOR4_X1 _11816_ ( .A1(_00889_ ), .A2(fanout_net_2 ), .A3(_04463_ ), .A4(_02459_ ), .ZN(_00254_ ) );
BUF_X4 _11817_ ( .A(_00855_ ), .Z(_04466_ ) );
NOR4_X1 _11818_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04463_ ), .A4(_02559_ ), .ZN(_00255_ ) );
AND3_X1 _11819_ ( .A1(_04465_ ), .A2(\de_pc [3] ), .A3(_04464_ ), .ZN(_00256_ ) );
NOR4_X1 _11820_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04463_ ), .A4(_02676_ ), .ZN(_00257_ ) );
NOR4_X1 _11821_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04463_ ), .A4(_02717_ ), .ZN(_00258_ ) );
NOR4_X1 _11822_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04463_ ), .A4(_02768_ ), .ZN(_00259_ ) );
AND3_X1 _11823_ ( .A1(_04465_ ), .A2(\de_pc [0] ), .A3(_04464_ ), .ZN(_00260_ ) );
AND3_X1 _11824_ ( .A1(_04465_ ), .A2(\de_pc [27] ), .A3(_04464_ ), .ZN(_00261_ ) );
NOR4_X1 _11825_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04463_ ), .A4(_02899_ ), .ZN(_00262_ ) );
AND3_X1 _11826_ ( .A1(_04465_ ), .A2(\de_pc [25] ), .A3(_04464_ ), .ZN(_00263_ ) );
AND3_X1 _11827_ ( .A1(_04465_ ), .A2(\de_pc [24] ), .A3(_04464_ ), .ZN(_00264_ ) );
BUF_X4 _11828_ ( .A(_00858_ ), .Z(_04467_ ) );
NOR4_X1 _11829_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04467_ ), .A4(_03025_ ), .ZN(_00265_ ) );
CLKBUF_X2 _11830_ ( .A(_00865_ ), .Z(_04468_ ) );
AND3_X1 _11831_ ( .A1(_04465_ ), .A2(\de_pc [22] ), .A3(_04468_ ), .ZN(_00266_ ) );
NAND4_X1 _11832_ ( .A1(_00750_ ), .A2(_00729_ ), .A3(_00728_ ), .A4(_00867_ ), .ZN(_04469_ ) );
NOR4_X1 _11833_ ( .A1(flush_$_OR__Y_B ), .A2(_00882_ ), .A3(_00705_ ), .A4(_04469_ ), .ZN(_00267_ ) );
NOR4_X1 _11834_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04467_ ), .A4(_04469_ ), .ZN(_00268_ ) );
BUF_X4 _11835_ ( .A(_02455_ ), .Z(_04470_ ) );
NOR3_X1 _11836_ ( .A1(_03512_ ), .A2(_04470_ ), .A3(_03576_ ), .ZN(_00269_ ) );
NOR3_X1 _11837_ ( .A1(_03588_ ), .A2(_04470_ ), .A3(_03627_ ), .ZN(_00270_ ) );
NOR3_X1 _11838_ ( .A1(_03635_ ), .A2(_04470_ ), .A3(_03663_ ), .ZN(_00271_ ) );
NOR2_X1 _11839_ ( .A1(_03705_ ), .A2(_04461_ ), .ZN(_00272_ ) );
NOR2_X1 _11840_ ( .A1(_03735_ ), .A2(_04461_ ), .ZN(_00273_ ) );
BUF_X4 _11841_ ( .A(_02455_ ), .Z(_04471_ ) );
NOR2_X1 _11842_ ( .A1(_03764_ ), .A2(_04471_ ), .ZN(_00274_ ) );
NOR3_X1 _11843_ ( .A1(_03768_ ), .A2(_04470_ ), .A3(_03789_ ), .ZN(_00275_ ) );
NOR2_X1 _11844_ ( .A1(_03815_ ), .A2(_04471_ ), .ZN(_00276_ ) );
NOR2_X1 _11845_ ( .A1(_03838_ ), .A2(_04471_ ), .ZN(_00277_ ) );
NOR2_X1 _11846_ ( .A1(_03861_ ), .A2(_04471_ ), .ZN(_00278_ ) );
NOR2_X1 _11847_ ( .A1(_03888_ ), .A2(_04471_ ), .ZN(_00279_ ) );
NOR2_X1 _11848_ ( .A1(_03913_ ), .A2(_04471_ ), .ZN(_00280_ ) );
NOR2_X1 _11849_ ( .A1(_03941_ ), .A2(_04471_ ), .ZN(_00281_ ) );
NOR2_X1 _11850_ ( .A1(_03968_ ), .A2(_04471_ ), .ZN(_00282_ ) );
NOR2_X1 _11851_ ( .A1(_03993_ ), .A2(_04471_ ), .ZN(_00283_ ) );
NOR2_X1 _11852_ ( .A1(_04018_ ), .A2(_04471_ ), .ZN(_00284_ ) );
BUF_X4 _11853_ ( .A(_02455_ ), .Z(_04472_ ) );
NOR2_X1 _11854_ ( .A1(_04043_ ), .A2(_04472_ ), .ZN(_00285_ ) );
BUF_X4 _11855_ ( .A(_00891_ ), .Z(_04473_ ) );
BUF_X4 _11856_ ( .A(_04473_ ), .Z(_04474_ ) );
OAI211_X1 _11857_ ( .A(_04474_ ), .B(_04069_ ), .C1(\ar_data [7] ), .C2(_04070_ ), .ZN(_04475_ ) );
INV_X1 _11858_ ( .A(_04475_ ), .ZN(_00286_ ) );
BUF_X2 _11859_ ( .A(_04473_ ), .Z(_04476_ ) );
OAI211_X1 _11860_ ( .A(_04102_ ), .B(_04476_ ), .C1(\ar_data [6] ), .C2(_04070_ ), .ZN(_04477_ ) );
INV_X1 _11861_ ( .A(_04477_ ), .ZN(_00287_ ) );
OAI211_X1 _11862_ ( .A(_04474_ ), .B(_04126_ ), .C1(\ar_data [5] ), .C2(_04070_ ), .ZN(_04478_ ) );
INV_X1 _11863_ ( .A(_04478_ ), .ZN(_00288_ ) );
OAI211_X1 _11864_ ( .A(_04474_ ), .B(_04152_ ), .C1(\ar_data [4] ), .C2(_04070_ ), .ZN(_04479_ ) );
INV_X1 _11865_ ( .A(_04479_ ), .ZN(_00289_ ) );
OAI211_X1 _11866_ ( .A(_04474_ ), .B(_04180_ ), .C1(\ar_data [3] ), .C2(_04070_ ), .ZN(_04480_ ) );
INV_X1 _11867_ ( .A(_04480_ ), .ZN(_00290_ ) );
OAI211_X1 _11868_ ( .A(_04474_ ), .B(_04204_ ), .C1(\ar_data [2] ), .C2(_04070_ ), .ZN(_04481_ ) );
INV_X1 _11869_ ( .A(_04481_ ), .ZN(_00291_ ) );
NOR3_X1 _11870_ ( .A1(_04215_ ), .A2(_04470_ ), .A3(_04236_ ), .ZN(_00292_ ) );
OAI211_X1 _11871_ ( .A(_04474_ ), .B(_04265_ ), .C1(\ar_data [1] ), .C2(_04070_ ), .ZN(_04482_ ) );
INV_X1 _11872_ ( .A(_04482_ ), .ZN(_00293_ ) );
OR2_X1 _11873_ ( .A1(_04070_ ), .A2(\ar_data [0] ), .ZN(_04483_ ) );
AND4_X1 _11874_ ( .A1(_04476_ ), .A2(_04483_ ), .A3(_03516_ ), .A4(_04288_ ), .ZN(_00294_ ) );
NOR2_X1 _11875_ ( .A1(_04319_ ), .A2(_04472_ ), .ZN(_00295_ ) );
NOR3_X1 _11876_ ( .A1(_04326_ ), .A2(_04470_ ), .A3(_04349_ ), .ZN(_00296_ ) );
NOR2_X1 _11877_ ( .A1(_04377_ ), .A2(_04472_ ), .ZN(_00297_ ) );
AND4_X1 _11878_ ( .A1(_04476_ ), .A2(_04382_ ), .A3(_03516_ ), .A4(_04399_ ), .ZN(_00298_ ) );
NOR2_X1 _11879_ ( .A1(_04424_ ), .A2(_04472_ ), .ZN(_00299_ ) );
NOR2_X1 _11880_ ( .A1(_04450_ ), .A2(_04472_ ), .ZN(_00300_ ) );
INV_X1 _11881_ ( .A(\u_exu.exe_start ), .ZN(_04484_ ) );
NOR2_X1 _11882_ ( .A1(_04484_ ), .A2(exu_valid ), .ZN(\u_exu.exe_end_$_ANDNOT__B_Y ) );
INV_X1 _11883_ ( .A(\u_exu.exe_end_$_ANDNOT__B_Y ), .ZN(_04485_ ) );
NOR4_X1 _11884_ ( .A1(_04466_ ), .A2(fanout_net_2 ), .A3(_04467_ ), .A4(_04485_ ), .ZN(_00301_ ) );
CLKBUF_X2 _11885_ ( .A(_03400_ ), .Z(_04486_ ) );
CLKBUF_X2 _11886_ ( .A(_03490_ ), .Z(_04487_ ) );
AND4_X1 _11887_ ( .A1(_03395_ ), .A2(_04486_ ), .A3(_04487_ ), .A4(fanout_net_19 ), .ZN(_04488_ ) );
NOR2_X1 _11888_ ( .A1(_03395_ ), .A2(fanout_net_13 ), .ZN(_04489_ ) );
BUF_X2 _11889_ ( .A(_03470_ ), .Z(_04490_ ) );
BUF_X2 _11890_ ( .A(_04490_ ), .Z(_04491_ ) );
AND2_X1 _11891_ ( .A1(_04489_ ), .A2(_04491_ ), .ZN(_04492_ ) );
BUF_X2 _11892_ ( .A(_03099_ ), .Z(_04493_ ) );
BUF_X4 _11893_ ( .A(_03100_ ), .Z(_04494_ ) );
BUF_X2 _11894_ ( .A(_04494_ ), .Z(_04495_ ) );
NAND4_X1 _11895_ ( .A1(_04492_ ), .A2(_04493_ ), .A3(_04495_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B_$_MUX__B_A_$_NAND__Y_B ), .ZN(_04496_ ) );
INV_X1 _11896_ ( .A(\u_exu.alu_ctrl [1] ), .ZN(_04497_ ) );
MUX2_X1 _11897_ ( .A(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ), .B(_04496_ ), .S(_04497_ ), .Z(_04498_ ) );
NOR2_X1 _11898_ ( .A1(_04498_ ), .A2(_03437_ ), .ZN(_04499_ ) );
OAI211_X1 _11899_ ( .A(_03401_ ), .B(fanout_net_19 ), .C1(fanout_net_11 ), .C2(\u_exu.alu_p2 [31] ), .ZN(_04500_ ) );
NAND2_X1 _11900_ ( .A1(fanout_net_11 ), .A2(\u_exu.alu_p2 [31] ), .ZN(_04501_ ) );
AOI21_X1 _11901_ ( .A(_04500_ ), .B1(_03395_ ), .B2(_04501_ ), .ZN(_04502_ ) );
AND2_X1 _11902_ ( .A1(_03142_ ), .A2(_03482_ ), .ZN(_04503_ ) );
OR3_X1 _11903_ ( .A1(_04499_ ), .A2(_04502_ ), .A3(_04503_ ), .ZN(_04504_ ) );
AND2_X2 _11904_ ( .A1(_03104_ ), .A2(\u_exu.alu_p2 [4] ), .ZN(_04505_ ) );
BUF_X2 _11905_ ( .A(_04505_ ), .Z(_04506_ ) );
BUF_X2 _11906_ ( .A(_03099_ ), .Z(_04507_ ) );
BUF_X2 _11907_ ( .A(_04507_ ), .Z(_04508_ ) );
AND2_X1 _11908_ ( .A1(_03089_ ), .A2(\u_exu.alu_p1 [15] ), .ZN(_04509_ ) );
AND2_X1 _11909_ ( .A1(\u_exu.alu_p1 [14] ), .A2(fanout_net_13 ), .ZN(_04510_ ) );
OR3_X1 _11910_ ( .A1(_04509_ ), .A2(fanout_net_14 ), .A3(_04510_ ), .ZN(_04511_ ) );
AND2_X1 _11911_ ( .A1(\u_exu.alu_p1 [12] ), .A2(fanout_net_13 ), .ZN(_04512_ ) );
INV_X1 _11912_ ( .A(_04512_ ), .ZN(_04513_ ) );
OAI211_X1 _11913_ ( .A(_04513_ ), .B(fanout_net_14 ), .C1(_03231_ ), .C2(fanout_net_13 ), .ZN(_04514_ ) );
AOI21_X1 _11914_ ( .A(fanout_net_16 ), .B1(_04511_ ), .B2(_04514_ ), .ZN(_04515_ ) );
BUF_X2 _11915_ ( .A(_03102_ ), .Z(_04516_ ) );
AND2_X1 _11916_ ( .A1(_03089_ ), .A2(\u_exu.alu_p1 [9] ), .ZN(_04517_ ) );
AND2_X1 _11917_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [8] ), .ZN(_04518_ ) );
OR3_X1 _11918_ ( .A1(_04517_ ), .A2(_04490_ ), .A3(_04518_ ), .ZN(_04519_ ) );
AND2_X1 _11919_ ( .A1(_03089_ ), .A2(\u_exu.alu_p1 [11] ), .ZN(_04520_ ) );
INV_X1 _11920_ ( .A(_04520_ ), .ZN(_04521_ ) );
AND2_X1 _11921_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [10] ), .ZN(_04522_ ) );
INV_X1 _11922_ ( .A(_04522_ ), .ZN(_04523_ ) );
NAND3_X1 _11923_ ( .A1(_04521_ ), .A2(_04491_ ), .A3(_04523_ ), .ZN(_04524_ ) );
AOI21_X1 _11924_ ( .A(_04516_ ), .B1(_04519_ ), .B2(_04524_ ), .ZN(_04525_ ) );
OAI21_X1 _11925_ ( .A(_04508_ ), .B1(_04515_ ), .B2(_04525_ ), .ZN(_04526_ ) );
BUF_X2 _11926_ ( .A(_03470_ ), .Z(_04527_ ) );
BUF_X2 _11927_ ( .A(_04527_ ), .Z(_04528_ ) );
AND2_X1 _11928_ ( .A1(_03089_ ), .A2(\u_exu.alu_p1 [7] ), .ZN(_04529_ ) );
AND2_X1 _11929_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [6] ), .ZN(_04530_ ) );
OAI21_X1 _11930_ ( .A(_04528_ ), .B1(_04529_ ), .B2(_04530_ ), .ZN(_04531_ ) );
AND2_X1 _11931_ ( .A1(_03088_ ), .A2(\u_exu.alu_p1 [5] ), .ZN(_04532_ ) );
AND2_X1 _11932_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [4] ), .ZN(_04533_ ) );
OAI21_X1 _11933_ ( .A(fanout_net_14 ), .B1(_04532_ ), .B2(_04533_ ), .ZN(_04534_ ) );
NAND2_X1 _11934_ ( .A1(_04531_ ), .A2(_04534_ ), .ZN(_04535_ ) );
NAND2_X1 _11935_ ( .A1(_04535_ ), .A2(_04516_ ), .ZN(_04536_ ) );
BUF_X2 _11936_ ( .A(_04494_ ), .Z(_04537_ ) );
BUF_X2 _11937_ ( .A(_04537_ ), .Z(_04538_ ) );
AND2_X1 _11938_ ( .A1(_03089_ ), .A2(\u_exu.alu_p1 [3] ), .ZN(_04539_ ) );
AND2_X1 _11939_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [2] ), .ZN(_04540_ ) );
OR3_X1 _11940_ ( .A1(_04539_ ), .A2(fanout_net_14 ), .A3(_04540_ ), .ZN(_04541_ ) );
INV_X1 _11941_ ( .A(\u_exu.alu_p1 [1] ), .ZN(_04542_ ) );
OAI211_X1 _11942_ ( .A(_03486_ ), .B(fanout_net_14 ), .C1(fanout_net_13 ), .C2(_04542_ ), .ZN(_04543_ ) );
NAND2_X1 _11943_ ( .A1(_04541_ ), .A2(_04543_ ), .ZN(_04544_ ) );
OAI211_X1 _11944_ ( .A(_04536_ ), .B(fanout_net_18 ), .C1(_04538_ ), .C2(_04544_ ), .ZN(_04545_ ) );
AND2_X1 _11945_ ( .A1(_04526_ ), .A2(_04545_ ), .ZN(_04546_ ) );
XNOR2_X1 _11946_ ( .A(_03394_ ), .B(_03396_ ), .ZN(_04547_ ) );
AND2_X1 _11947_ ( .A1(_03087_ ), .A2(fanout_net_19 ), .ZN(_04548_ ) );
BUF_X2 _11948_ ( .A(_04548_ ), .Z(_04549_ ) );
BUF_X4 _11949_ ( .A(_04549_ ), .Z(_04550_ ) );
AOI221_X2 _11950_ ( .A(_04504_ ), .B1(_04506_ ), .B2(_04546_ ), .C1(_04547_ ), .C2(_04550_ ), .ZN(_04551_ ) );
NOR2_X1 _11951_ ( .A1(_03177_ ), .A2(fanout_net_13 ), .ZN(_04552_ ) );
AND2_X1 _11952_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [28] ), .ZN(_04553_ ) );
NOR2_X1 _11953_ ( .A1(_04552_ ), .A2(_04553_ ), .ZN(_04554_ ) );
NOR2_X1 _11954_ ( .A1(_04554_ ), .A2(_04491_ ), .ZN(_04555_ ) );
AND3_X1 _11955_ ( .A1(_04491_ ), .A2(\u_exu.alu_p1 [30] ), .A3(fanout_net_13 ), .ZN(_04556_ ) );
OR4_X1 _11956_ ( .A1(fanout_net_16 ), .A2(_04555_ ), .A3(_04492_ ), .A4(_04556_ ), .ZN(_04557_ ) );
AND2_X1 _11957_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [26] ), .ZN(_04558_ ) );
INV_X1 _11958_ ( .A(_04558_ ), .ZN(_04559_ ) );
OAI211_X1 _11959_ ( .A(_04559_ ), .B(_03470_ ), .C1(fanout_net_13 ), .C2(_03355_ ), .ZN(_04560_ ) );
NOR2_X1 _11960_ ( .A1(_03370_ ), .A2(fanout_net_13 ), .ZN(_04561_ ) );
INV_X1 _11961_ ( .A(_04561_ ), .ZN(_04562_ ) );
AND2_X1 _11962_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [24] ), .ZN(_04563_ ) );
INV_X1 _11963_ ( .A(_04563_ ), .ZN(_04564_ ) );
NAND3_X1 _11964_ ( .A1(_04562_ ), .A2(fanout_net_14 ), .A3(_04564_ ), .ZN(_04565_ ) );
AND2_X1 _11965_ ( .A1(_04560_ ), .A2(_04565_ ), .ZN(_04566_ ) );
OR2_X1 _11966_ ( .A1(_04566_ ), .A2(_04538_ ), .ZN(_04567_ ) );
AOI21_X1 _11967_ ( .A(fanout_net_18 ), .B1(_04557_ ), .B2(_04567_ ), .ZN(_04568_ ) );
AND2_X1 _11968_ ( .A1(_03089_ ), .A2(\u_exu.alu_p1 [17] ), .ZN(_04569_ ) );
AND2_X1 _11969_ ( .A1(\u_exu.alu_p1 [16] ), .A2(fanout_net_13 ), .ZN(_04570_ ) );
OR3_X1 _11970_ ( .A1(_04569_ ), .A2(_04527_ ), .A3(_04570_ ), .ZN(_04571_ ) );
AND2_X1 _11971_ ( .A1(_03089_ ), .A2(\u_exu.alu_p1 [19] ), .ZN(_04572_ ) );
AND2_X1 _11972_ ( .A1(\u_exu.alu_p1 [18] ), .A2(fanout_net_13 ), .ZN(_04573_ ) );
OR3_X1 _11973_ ( .A1(_04572_ ), .A2(fanout_net_14 ), .A3(_04573_ ), .ZN(_04574_ ) );
NAND3_X1 _11974_ ( .A1(_04571_ ), .A2(_04574_ ), .A3(fanout_net_16 ), .ZN(_04575_ ) );
AND2_X1 _11975_ ( .A1(_03088_ ), .A2(\u_exu.alu_p1 [21] ), .ZN(_04576_ ) );
INV_X1 _11976_ ( .A(_04576_ ), .ZN(_04577_ ) );
AND2_X1 _11977_ ( .A1(\u_exu.alu_p1 [20] ), .A2(fanout_net_13 ), .ZN(_04578_ ) );
INV_X1 _11978_ ( .A(_04578_ ), .ZN(_04579_ ) );
NAND3_X1 _11979_ ( .A1(_04577_ ), .A2(fanout_net_14 ), .A3(_04579_ ), .ZN(_04580_ ) );
NOR2_X1 _11980_ ( .A1(_03295_ ), .A2(fanout_net_13 ), .ZN(_04581_ ) );
INV_X1 _11981_ ( .A(_04581_ ), .ZN(_04582_ ) );
AND2_X1 _11982_ ( .A1(fanout_net_13 ), .A2(\u_exu.alu_p1 [22] ), .ZN(_04583_ ) );
INV_X1 _11983_ ( .A(_04583_ ), .ZN(_04584_ ) );
NAND3_X1 _11984_ ( .A1(_04582_ ), .A2(_03470_ ), .A3(_04584_ ), .ZN(_04585_ ) );
NAND3_X1 _11985_ ( .A1(_04580_ ), .A2(_04516_ ), .A3(_04585_ ), .ZN(_04586_ ) );
AND3_X1 _11986_ ( .A1(_04575_ ), .A2(fanout_net_18 ), .A3(_04586_ ), .ZN(_04587_ ) );
AND2_X1 _11987_ ( .A1(_03104_ ), .A2(_03098_ ), .ZN(_04588_ ) );
INV_X1 _11988_ ( .A(_04588_ ), .ZN(_04589_ ) );
NOR3_X1 _11989_ ( .A1(_04568_ ), .A2(_04587_ ), .A3(_04589_ ), .ZN(_04590_ ) );
NOR2_X1 _11990_ ( .A1(_04590_ ), .A2(_03079_ ), .ZN(_04591_ ) );
AOI21_X1 _11991_ ( .A(_04488_ ), .B1(_04551_ ), .B2(_04591_ ), .ZN(_04592_ ) );
CLKBUF_X2 _11992_ ( .A(_04473_ ), .Z(_04593_ ) );
NAND2_X1 _11993_ ( .A1(_04592_ ), .A2(_04593_ ), .ZN(_04594_ ) );
INV_X1 _11994_ ( .A(_04594_ ), .ZN(_00303_ ) );
NOR2_X1 _11995_ ( .A1(_01113_ ), .A2(_00700_ ), .ZN(_04595_ ) );
NAND2_X1 _11996_ ( .A1(_04595_ ), .A2(_00704_ ), .ZN(_04596_ ) );
AOI211_X1 _11997_ ( .A(_00894_ ), .B(_04485_ ), .C1(_00746_ ), .C2(_04596_ ), .ZN(_00304_ ) );
XNOR2_X1 _11998_ ( .A(_03387_ ), .B(_03390_ ), .ZN(_04597_ ) );
AND2_X1 _11999_ ( .A1(_04597_ ), .A2(_04549_ ), .ZN(_04598_ ) );
NOR2_X1 _12000_ ( .A1(_04497_ ), .A2(\u_exu.alu_p2 [4] ), .ZN(_04599_ ) );
OR3_X1 _12001_ ( .A1(_03460_ ), .A2(fanout_net_16 ), .A3(fanout_net_14 ), .ZN(_04600_ ) );
OAI21_X1 _12002_ ( .A(\u_exu.alu_p1 [31] ), .B1(fanout_net_16 ), .B2(fanout_net_14 ), .ZN(_04601_ ) );
AOI21_X1 _12003_ ( .A(fanout_net_18 ), .B1(_04600_ ), .B2(_04601_ ), .ZN(_04602_ ) );
AND2_X1 _12004_ ( .A1(\u_exu.alu_p1 [31] ), .A2(fanout_net_18 ), .ZN(_04603_ ) );
OAI21_X1 _12005_ ( .A(_04599_ ), .B1(_04602_ ), .B2(_04603_ ), .ZN(_04604_ ) );
AND2_X1 _12006_ ( .A1(\u_exu.alu_ctrl [1] ), .A2(\u_exu.alu_p2 [4] ), .ZN(_04605_ ) );
AND2_X1 _12007_ ( .A1(_04605_ ), .A2(\u_exu.alu_p1 [31] ), .ZN(_04606_ ) );
NOR2_X1 _12008_ ( .A1(_04600_ ), .A2(fanout_net_18 ), .ZN(_04607_ ) );
NOR2_X1 _12009_ ( .A1(\u_exu.alu_ctrl [1] ), .A2(\u_exu.alu_p2 [4] ), .ZN(_04608_ ) );
AOI21_X1 _12010_ ( .A(_04606_ ), .B1(_04607_ ), .B2(_04608_ ), .ZN(_04609_ ) );
AOI21_X1 _12011_ ( .A(_03437_ ), .B1(_04604_ ), .B2(_04609_ ), .ZN(_04610_ ) );
OAI211_X1 _12012_ ( .A(_03466_ ), .B(fanout_net_14 ), .C1(fanout_net_13 ), .C2(_03182_ ), .ZN(_04611_ ) );
MUX2_X1 _12013_ ( .A(\u_exu.alu_p1 [30] ), .B(\u_exu.alu_p1 [29] ), .S(\u_exu.alu_p2 [0] ), .Z(_04612_ ) );
OAI211_X1 _12014_ ( .A(_04611_ ), .B(_04495_ ), .C1(fanout_net_14 ), .C2(_04612_ ), .ZN(_04613_ ) );
NOR2_X1 _12015_ ( .A1(_03463_ ), .A2(_03471_ ), .ZN(_04614_ ) );
NOR2_X1 _12016_ ( .A1(_03468_ ), .A2(_03451_ ), .ZN(_04615_ ) );
MUX2_X1 _12017_ ( .A(_04614_ ), .B(_04615_ ), .S(fanout_net_14 ), .Z(_04616_ ) );
OAI211_X1 _12018_ ( .A(_04613_ ), .B(_04507_ ), .C1(_04616_ ), .C2(_04516_ ), .ZN(_04617_ ) );
BUF_X2 _12019_ ( .A(_03098_ ), .Z(_04618_ ) );
OR3_X1 _12020_ ( .A1(_03448_ ), .A2(_03441_ ), .A3(_04528_ ), .ZN(_04619_ ) );
NOR2_X1 _12021_ ( .A1(_03299_ ), .A2(\u_exu.alu_p2 [0] ), .ZN(_04620_ ) );
OR3_X1 _12022_ ( .A1(_04620_ ), .A2(_03449_ ), .A3(fanout_net_14 ), .ZN(_04621_ ) );
NAND3_X1 _12023_ ( .A1(_04619_ ), .A2(_04621_ ), .A3(_04537_ ), .ZN(_04622_ ) );
OR3_X1 _12024_ ( .A1(_03443_ ), .A2(_03427_ ), .A3(_04528_ ), .ZN(_04623_ ) );
OR3_X1 _12025_ ( .A1(_03440_ ), .A2(_03444_ ), .A3(fanout_net_14 ), .ZN(_04624_ ) );
NAND3_X1 _12026_ ( .A1(_04623_ ), .A2(_04624_ ), .A3(fanout_net_16 ), .ZN(_04625_ ) );
NAND3_X1 _12027_ ( .A1(_04622_ ), .A2(_04625_ ), .A3(fanout_net_18 ), .ZN(_04626_ ) );
AND3_X1 _12028_ ( .A1(_04617_ ), .A2(_04618_ ), .A3(_04626_ ), .ZN(_04627_ ) );
AND3_X1 _12029_ ( .A1(_04627_ ), .A2(\u_exu.alu_ctrl [6] ), .A3(_03078_ ), .ZN(_04628_ ) );
BUF_X4 _12030_ ( .A(_03099_ ), .Z(_04629_ ) );
BUF_X4 _12031_ ( .A(_04629_ ), .Z(_04630_ ) );
OR3_X1 _12032_ ( .A1(_03422_ ), .A2(_03415_ ), .A3(_04528_ ), .ZN(_04631_ ) );
OR3_X1 _12033_ ( .A1(_03419_ ), .A2(_03423_ ), .A3(fanout_net_14 ), .ZN(_04632_ ) );
AOI21_X1 _12034_ ( .A(_04537_ ), .B1(_04631_ ), .B2(_04632_ ), .ZN(_04633_ ) );
OAI21_X1 _12035_ ( .A(_04491_ ), .B1(_03426_ ), .B2(_03430_ ), .ZN(_04634_ ) );
OAI21_X1 _12036_ ( .A(fanout_net_14 ), .B1(_03429_ ), .B2(_03420_ ), .ZN(_04635_ ) );
AND3_X1 _12037_ ( .A1(_04634_ ), .A2(_04635_ ), .A3(_04495_ ), .ZN(_04636_ ) );
OAI21_X1 _12038_ ( .A(_04630_ ), .B1(_04633_ ), .B2(_04636_ ), .ZN(_04637_ ) );
OR3_X1 _12039_ ( .A1(_03411_ ), .A2(_03406_ ), .A3(_04490_ ), .ZN(_04638_ ) );
OR3_X1 _12040_ ( .A1(_03414_ ), .A2(_03412_ ), .A3(fanout_net_14 ), .ZN(_04639_ ) );
NAND3_X1 _12041_ ( .A1(_04638_ ), .A2(_04639_ ), .A3(_03102_ ), .ZN(_04640_ ) );
AND2_X1 _12042_ ( .A1(\u_exu.alu_p2 [0] ), .A2(\u_exu.alu_p1 [1] ), .ZN(_04641_ ) );
OR3_X1 _12043_ ( .A1(_03405_ ), .A2(_04641_ ), .A3(fanout_net_14 ), .ZN(_04642_ ) );
OAI21_X1 _12044_ ( .A(_04642_ ), .B1(_04491_ ), .B2(_03095_ ), .ZN(_04643_ ) );
OAI211_X1 _12045_ ( .A(_04640_ ), .B(fanout_net_18 ), .C1(_04643_ ), .C2(_04538_ ), .ZN(_04644_ ) );
NAND3_X1 _12046_ ( .A1(_04637_ ), .A2(_04644_ ), .A3(_04506_ ), .ZN(_04645_ ) );
BUF_X2 _12047_ ( .A(_03482_ ), .Z(_04646_ ) );
NAND2_X1 _12048_ ( .A1(_03121_ ), .A2(_04646_ ), .ZN(_04647_ ) );
AOI21_X1 _12049_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [30] ), .B2(\u_exu.alu_p2 [30] ), .ZN(_04648_ ) );
BUF_X4 _12050_ ( .A(_03401_ ), .Z(_04649_ ) );
OAI211_X1 _12051_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [30] ), .C2(\u_exu.alu_p2 [30] ), .ZN(_04650_ ) );
OAI211_X1 _12052_ ( .A(_04645_ ), .B(_04647_ ), .C1(_04648_ ), .C2(_04650_ ), .ZN(_04651_ ) );
NOR4_X1 _12053_ ( .A1(_04598_ ), .A2(_04610_ ), .A3(_04628_ ), .A4(_04651_ ), .ZN(_04652_ ) );
BUF_X4 _12054_ ( .A(_03080_ ), .Z(_04653_ ) );
MUX2_X1 _12055_ ( .A(_03389_ ), .B(_04652_ ), .S(_04653_ ), .Z(_04654_ ) );
OR2_X1 _12056_ ( .A1(_04654_ ), .A2(_02455_ ), .ZN(_04655_ ) );
INV_X1 _12057_ ( .A(_04655_ ), .ZN(_00305_ ) );
NAND2_X1 _12058_ ( .A1(_03292_ ), .A2(_03326_ ), .ZN(_04656_ ) );
AND2_X2 _12059_ ( .A1(_04656_ ), .A2(_03339_ ), .ZN(_04657_ ) );
NOR2_X1 _12060_ ( .A1(_03303_ ), .A2(\u_exu.alu_p1 [20] ), .ZN(_04658_ ) );
NOR3_X1 _12061_ ( .A1(_04657_ ), .A2(_03342_ ), .A3(_04658_ ), .ZN(_04659_ ) );
OR3_X2 _12062_ ( .A1(_04659_ ), .A2(_03308_ ), .A3(_03342_ ), .ZN(_04660_ ) );
OAI21_X1 _12063_ ( .A(_03308_ ), .B1(_04659_ ), .B2(_03342_ ), .ZN(_04661_ ) );
AND3_X2 _12064_ ( .A1(_04660_ ), .A2(_04548_ ), .A3(_04661_ ), .ZN(_04662_ ) );
NAND3_X1 _12065_ ( .A1(_04577_ ), .A2(_03470_ ), .A3(_04584_ ), .ZN(_04663_ ) );
NAND3_X1 _12066_ ( .A1(_04582_ ), .A2(fanout_net_15 ), .A3(_04564_ ), .ZN(_04664_ ) );
AOI21_X1 _12067_ ( .A(fanout_net_16 ), .B1(_04663_ ), .B2(_04664_ ), .ZN(_04665_ ) );
NOR2_X1 _12068_ ( .A1(_04561_ ), .A2(_04558_ ), .ZN(_04666_ ) );
NOR2_X1 _12069_ ( .A1(_03355_ ), .A2(\u_exu.alu_p2 [0] ), .ZN(_04667_ ) );
NOR2_X1 _12070_ ( .A1(_04667_ ), .A2(_04553_ ), .ZN(_04668_ ) );
MUX2_X1 _12071_ ( .A(_04666_ ), .B(_04668_ ), .S(fanout_net_15 ), .Z(_04669_ ) );
AOI21_X1 _12072_ ( .A(_04665_ ), .B1(fanout_net_16 ), .B2(_04669_ ), .ZN(_04670_ ) );
AND2_X1 _12073_ ( .A1(_04670_ ), .A2(_03099_ ), .ZN(_04671_ ) );
INV_X1 _12074_ ( .A(_04489_ ), .ZN(_04672_ ) );
MUX2_X1 _12075_ ( .A(_03177_ ), .B(_03389_ ), .S(\u_exu.alu_p2 [0] ), .Z(_04673_ ) );
MUX2_X1 _12076_ ( .A(_04672_ ), .B(_04673_ ), .S(_03470_ ), .Z(_04674_ ) );
NOR3_X1 _12077_ ( .A1(_04674_ ), .A2(_03099_ ), .A3(fanout_net_16 ), .ZN(_04675_ ) );
OAI21_X1 _12078_ ( .A(_04608_ ), .B1(_04671_ ), .B2(_04675_ ), .ZN(_04676_ ) );
INV_X1 _12079_ ( .A(_04606_ ), .ZN(_04677_ ) );
AND2_X1 _12080_ ( .A1(\u_exu.alu_p1 [31] ), .A2(fanout_net_16 ), .ZN(_04678_ ) );
INV_X1 _12081_ ( .A(_04678_ ), .ZN(_04679_ ) );
MUX2_X1 _12082_ ( .A(_03395_ ), .B(_04673_ ), .S(_03096_ ), .Z(_04680_ ) );
OAI21_X1 _12083_ ( .A(_04679_ ), .B1(_04680_ ), .B2(fanout_net_16 ), .ZN(_04681_ ) );
AND2_X1 _12084_ ( .A1(_04681_ ), .A2(fanout_net_18 ), .ZN(_04682_ ) );
NOR2_X1 _12085_ ( .A1(_04671_ ), .A2(_04682_ ), .ZN(_04683_ ) );
INV_X1 _12086_ ( .A(_04599_ ), .ZN(_04684_ ) );
OAI211_X1 _12087_ ( .A(_04676_ ), .B(_04677_ ), .C1(_04683_ ), .C2(_04684_ ), .ZN(_04685_ ) );
BUF_X4 _12088_ ( .A(_03436_ ), .Z(_04686_ ) );
AND2_X1 _12089_ ( .A1(_04685_ ), .A2(_04686_ ), .ZN(_04687_ ) );
OAI21_X1 _12090_ ( .A(_04490_ ), .B1(_04576_ ), .B2(_04578_ ), .ZN(_04688_ ) );
OAI21_X1 _12091_ ( .A(fanout_net_15 ), .B1(_04572_ ), .B2(_04573_ ), .ZN(_04689_ ) );
NAND2_X1 _12092_ ( .A1(_04688_ ), .A2(_04689_ ), .ZN(_04690_ ) );
NAND2_X1 _12093_ ( .A1(_04690_ ), .A2(_04494_ ), .ZN(_04691_ ) );
OAI21_X1 _12094_ ( .A(_04527_ ), .B1(_04569_ ), .B2(_04570_ ), .ZN(_04692_ ) );
OAI21_X1 _12095_ ( .A(fanout_net_15 ), .B1(_04509_ ), .B2(_04510_ ), .ZN(_04693_ ) );
NAND2_X1 _12096_ ( .A1(_04692_ ), .A2(_04693_ ), .ZN(_04694_ ) );
NAND2_X1 _12097_ ( .A1(_04694_ ), .A2(fanout_net_16 ), .ZN(_04695_ ) );
AOI21_X1 _12098_ ( .A(fanout_net_18 ), .B1(_04691_ ), .B2(_04695_ ), .ZN(_04696_ ) );
OAI21_X1 _12099_ ( .A(_04490_ ), .B1(_04517_ ), .B2(_04518_ ), .ZN(_04697_ ) );
OAI21_X1 _12100_ ( .A(fanout_net_15 ), .B1(_04529_ ), .B2(_04530_ ), .ZN(_04698_ ) );
NAND2_X1 _12101_ ( .A1(_04697_ ), .A2(_04698_ ), .ZN(_04699_ ) );
NAND2_X1 _12102_ ( .A1(_04699_ ), .A2(fanout_net_16 ), .ZN(_04700_ ) );
OAI21_X1 _12103_ ( .A(fanout_net_15 ), .B1(_04520_ ), .B2(_04522_ ), .ZN(_04701_ ) );
NOR2_X1 _12104_ ( .A1(_03231_ ), .A2(\u_exu.alu_p2 [0] ), .ZN(_04702_ ) );
OAI21_X1 _12105_ ( .A(_04490_ ), .B1(_04702_ ), .B2(_04512_ ), .ZN(_04703_ ) );
NAND2_X1 _12106_ ( .A1(_04701_ ), .A2(_04703_ ), .ZN(_04704_ ) );
NAND2_X1 _12107_ ( .A1(_04704_ ), .A2(_03102_ ), .ZN(_04705_ ) );
NAND2_X1 _12108_ ( .A1(_04700_ ), .A2(_04705_ ), .ZN(_04706_ ) );
AOI21_X1 _12109_ ( .A(_04696_ ), .B1(fanout_net_18 ), .B2(_04706_ ), .ZN(_04707_ ) );
NOR2_X1 _12110_ ( .A1(_04707_ ), .A2(_04589_ ), .ZN(_04708_ ) );
MUX2_X1 _12111_ ( .A(_04542_ ), .B(_03094_ ), .S(\u_exu.alu_p2 [0] ), .Z(_04709_ ) );
NOR2_X1 _12112_ ( .A1(_04709_ ), .A2(fanout_net_15 ), .ZN(_04710_ ) );
OAI21_X1 _12113_ ( .A(_03470_ ), .B1(_04532_ ), .B2(_04533_ ), .ZN(_04711_ ) );
OAI21_X1 _12114_ ( .A(fanout_net_15 ), .B1(_04539_ ), .B2(_04540_ ), .ZN(_04712_ ) );
NAND2_X1 _12115_ ( .A1(_04711_ ), .A2(_04712_ ), .ZN(_04713_ ) );
MUX2_X1 _12116_ ( .A(_04710_ ), .B(_04713_ ), .S(_03101_ ), .Z(_04714_ ) );
NAND3_X1 _12117_ ( .A1(_04714_ ), .A2(_04629_ ), .A3(_04505_ ), .ZN(_04715_ ) );
NAND2_X1 _12118_ ( .A1(_03114_ ), .A2(_03482_ ), .ZN(_04716_ ) );
AOI21_X1 _12119_ ( .A(\u_exu.alu_p1 [21] ), .B1(\u_exu.alu_p2 [21] ), .B2(fanout_net_11 ), .ZN(_04717_ ) );
OAI211_X1 _12120_ ( .A(_03401_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p2 [21] ), .C2(fanout_net_11 ), .ZN(_04718_ ) );
OAI211_X1 _12121_ ( .A(_04715_ ), .B(_04716_ ), .C1(_04717_ ), .C2(_04718_ ), .ZN(_04719_ ) );
OR4_X4 _12122_ ( .A1(_04662_ ), .A2(_04687_ ), .A3(_04708_ ), .A4(_04719_ ), .ZN(_04720_ ) );
MUX2_X2 _12123_ ( .A(\u_exu.alu_p1 [21] ), .B(_04720_ ), .S(_04653_ ), .Z(_04721_ ) );
AND2_X1 _12124_ ( .A1(_04721_ ), .A2(_04593_ ), .ZN(_00306_ ) );
AND4_X1 _12125_ ( .A1(_03304_ ), .A2(_04486_ ), .A3(_04487_ ), .A4(fanout_net_19 ), .ZN(_04722_ ) );
BUF_X4 _12126_ ( .A(_03435_ ), .Z(_04723_ ) );
BUF_X4 _12127_ ( .A(_04723_ ), .Z(_04724_ ) );
NOR4_X1 _12128_ ( .A1(_04659_ ), .A2(_04724_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_04487_ ), .ZN(_04725_ ) );
INV_X1 _12129_ ( .A(_04657_ ), .ZN(_04726_ ) );
OAI21_X1 _12130_ ( .A(_04725_ ), .B1(_03305_ ), .B2(_04726_ ), .ZN(_04727_ ) );
MUX2_X1 _12131_ ( .A(_03474_ ), .B(_03454_ ), .S(_03101_ ), .Z(_04728_ ) );
NOR2_X1 _12132_ ( .A1(_04728_ ), .A2(fanout_net_18 ), .ZN(_04729_ ) );
NOR3_X1 _12133_ ( .A1(_03461_ ), .A2(_04493_ ), .A3(fanout_net_16 ), .ZN(_04730_ ) );
NOR2_X1 _12134_ ( .A1(_04729_ ), .A2(_04730_ ), .ZN(_04731_ ) );
INV_X1 _12135_ ( .A(_04608_ ), .ZN(_04732_ ) );
OAI21_X1 _12136_ ( .A(_04679_ ), .B1(_03461_ ), .B2(fanout_net_16 ), .ZN(_04733_ ) );
AND2_X1 _12137_ ( .A1(_04733_ ), .A2(fanout_net_18 ), .ZN(_04734_ ) );
NOR2_X1 _12138_ ( .A1(_04729_ ), .A2(_04734_ ), .ZN(_04735_ ) );
OAI221_X1 _12139_ ( .A(_04677_ ), .B1(_04731_ ), .B2(_04732_ ), .C1(_04684_ ), .C2(_04735_ ), .ZN(_04736_ ) );
BUF_X4 _12140_ ( .A(_04686_ ), .Z(_04737_ ) );
NAND2_X1 _12141_ ( .A1(_04736_ ), .A2(_04737_ ), .ZN(_04738_ ) );
OAI21_X1 _12142_ ( .A(_04528_ ), .B1(_03422_ ), .B2(_03415_ ), .ZN(_04739_ ) );
OAI21_X1 _12143_ ( .A(fanout_net_15 ), .B1(_03414_ ), .B2(_03412_ ), .ZN(_04740_ ) );
NAND2_X1 _12144_ ( .A1(_04739_ ), .A2(_04740_ ), .ZN(_04741_ ) );
NAND2_X1 _12145_ ( .A1(_04741_ ), .A2(fanout_net_16 ), .ZN(_04742_ ) );
OR3_X1 _12146_ ( .A1(_03419_ ), .A2(_03423_ ), .A3(_04490_ ), .ZN(_04743_ ) );
OR3_X1 _12147_ ( .A1(_03429_ ), .A2(_03420_ ), .A3(fanout_net_15 ), .ZN(_04744_ ) );
NAND3_X1 _12148_ ( .A1(_04743_ ), .A2(_04744_ ), .A3(_04495_ ), .ZN(_04745_ ) );
NAND3_X1 _12149_ ( .A1(_04742_ ), .A2(_04745_ ), .A3(fanout_net_18 ), .ZN(_04746_ ) );
OAI21_X1 _12150_ ( .A(_04528_ ), .B1(_03443_ ), .B2(_03427_ ), .ZN(_04747_ ) );
OAI21_X1 _12151_ ( .A(fanout_net_15 ), .B1(_03426_ ), .B2(_03430_ ), .ZN(_04748_ ) );
NAND2_X1 _12152_ ( .A1(_04747_ ), .A2(_04748_ ), .ZN(_04749_ ) );
NAND2_X1 _12153_ ( .A1(_04749_ ), .A2(fanout_net_16 ), .ZN(_04750_ ) );
OR3_X1 _12154_ ( .A1(_03440_ ), .A2(_03444_ ), .A3(_04490_ ), .ZN(_04751_ ) );
OR3_X1 _12155_ ( .A1(_03448_ ), .A2(_03441_ ), .A3(fanout_net_15 ), .ZN(_04752_ ) );
NAND3_X1 _12156_ ( .A1(_04751_ ), .A2(_04752_ ), .A3(_04495_ ), .ZN(_04753_ ) );
BUF_X4 _12157_ ( .A(_04630_ ), .Z(_04754_ ) );
NAND3_X1 _12158_ ( .A1(_04750_ ), .A2(_04753_ ), .A3(_04754_ ), .ZN(_04755_ ) );
BUF_X2 _12159_ ( .A(_04588_ ), .Z(_04756_ ) );
BUF_X2 _12160_ ( .A(_04756_ ), .Z(_04757_ ) );
NAND3_X1 _12161_ ( .A1(_04746_ ), .A2(_04755_ ), .A3(_04757_ ), .ZN(_04758_ ) );
OAI21_X1 _12162_ ( .A(_04527_ ), .B1(_03411_ ), .B2(_03406_ ), .ZN(_04759_ ) );
OAI21_X1 _12163_ ( .A(fanout_net_15 ), .B1(_03405_ ), .B2(_04641_ ), .ZN(_04760_ ) );
NAND2_X1 _12164_ ( .A1(_04759_ ), .A2(_04760_ ), .ZN(_04761_ ) );
MUX2_X1 _12165_ ( .A(_03097_ ), .B(_04761_ ), .S(_03101_ ), .Z(_04762_ ) );
NAND3_X1 _12166_ ( .A1(_04762_ ), .A2(_04754_ ), .A3(_04506_ ), .ZN(_04763_ ) );
OAI211_X1 _12167_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [20] ), .C2(\u_exu.alu_p2 [20] ), .ZN(_04764_ ) );
AOI21_X1 _12168_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [20] ), .B2(\u_exu.alu_p2 [20] ), .ZN(_04765_ ) );
NOR2_X1 _12169_ ( .A1(_04764_ ), .A2(_04765_ ), .ZN(_04766_ ) );
BUF_X4 _12170_ ( .A(_03482_ ), .Z(_04767_ ) );
AOI211_X1 _12171_ ( .A(_03079_ ), .B(_04766_ ), .C1(_03155_ ), .C2(_04767_ ), .ZN(_04768_ ) );
AND4_X1 _12172_ ( .A1(_04738_ ), .A2(_04758_ ), .A3(_04763_ ), .A4(_04768_ ), .ZN(_04769_ ) );
AOI211_X1 _12173_ ( .A(_04460_ ), .B(_04722_ ), .C1(_04727_ ), .C2(_04769_ ), .ZN(_00307_ ) );
NOR4_X1 _12174_ ( .A1(_04724_ ), .A2(\u_exu.alu_p1 [19] ), .A3(\u_exu.alu_ctrl [5] ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_04770_ ) );
NAND2_X1 _12175_ ( .A1(_03292_ ), .A2(_03318_ ), .ZN(_04771_ ) );
AOI21_X1 _12176_ ( .A(_03332_ ), .B1(_04771_ ), .B2(_03331_ ), .ZN(_04772_ ) );
OR3_X1 _12177_ ( .A1(_04772_ ), .A2(_03321_ ), .A3(_03337_ ), .ZN(_04773_ ) );
OAI21_X1 _12178_ ( .A(_03321_ ), .B1(_04772_ ), .B2(_03337_ ), .ZN(_04774_ ) );
AND3_X1 _12179_ ( .A1(_04773_ ), .A2(_04549_ ), .A3(_04774_ ), .ZN(_04775_ ) );
NAND4_X1 _12180_ ( .A1(_04528_ ), .A2(_03089_ ), .A3(\u_exu.alu_p1 [31] ), .A4(fanout_net_16 ), .ZN(_04776_ ) );
MUX2_X1 _12181_ ( .A(_04668_ ), .B(_04673_ ), .S(fanout_net_15 ), .Z(_04777_ ) );
OAI21_X1 _12182_ ( .A(_04776_ ), .B1(_04777_ ), .B2(fanout_net_16 ), .ZN(_04778_ ) );
AND2_X1 _12183_ ( .A1(_04778_ ), .A2(fanout_net_18 ), .ZN(_04779_ ) );
OR3_X1 _12184_ ( .A1(_04572_ ), .A2(fanout_net_15 ), .A3(_04578_ ), .ZN(_04780_ ) );
NAND3_X1 _12185_ ( .A1(_04577_ ), .A2(fanout_net_15 ), .A3(_04584_ ), .ZN(_04781_ ) );
AOI21_X1 _12186_ ( .A(fanout_net_16 ), .B1(_04780_ ), .B2(_04781_ ), .ZN(_04782_ ) );
NAND3_X1 _12187_ ( .A1(_04562_ ), .A2(fanout_net_15 ), .A3(_04559_ ), .ZN(_04783_ ) );
NAND3_X1 _12188_ ( .A1(_04582_ ), .A2(_04490_ ), .A3(_04564_ ), .ZN(_04784_ ) );
AOI21_X1 _12189_ ( .A(_04494_ ), .B1(_04783_ ), .B2(_04784_ ), .ZN(_04785_ ) );
NOR3_X1 _12190_ ( .A1(_04782_ ), .A2(_04785_ ), .A3(fanout_net_18 ), .ZN(_04786_ ) );
OAI21_X1 _12191_ ( .A(_04608_ ), .B1(_04779_ ), .B2(_04786_ ), .ZN(_04787_ ) );
AND2_X1 _12192_ ( .A1(_04787_ ), .A2(_04677_ ), .ZN(_04788_ ) );
OR2_X1 _12193_ ( .A1(_04777_ ), .A2(fanout_net_16 ), .ZN(_04789_ ) );
AOI21_X1 _12194_ ( .A(_04629_ ), .B1(_04789_ ), .B2(_04679_ ), .ZN(_04790_ ) );
OAI21_X1 _12195_ ( .A(_04599_ ), .B1(_04790_ ), .B2(_04786_ ), .ZN(_04791_ ) );
AOI21_X1 _12196_ ( .A(_03437_ ), .B1(_04788_ ), .B2(_04791_ ), .ZN(_04792_ ) );
AND3_X1 _12197_ ( .A1(_04541_ ), .A2(_04516_ ), .A3(_04543_ ), .ZN(_04793_ ) );
AND3_X1 _12198_ ( .A1(_04793_ ), .A2(_04754_ ), .A3(_04506_ ), .ZN(_04794_ ) );
OR4_X1 _12199_ ( .A1(_03435_ ), .A2(_03151_ ), .A3(_03400_ ), .A4(_03490_ ), .ZN(_04795_ ) );
OAI211_X1 _12200_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(fanout_net_11 ), .C2(_03151_ ), .ZN(_04796_ ) );
AOI21_X1 _12201_ ( .A(_03150_ ), .B1(_04795_ ), .B2(_04796_ ), .ZN(_04797_ ) );
NOR4_X1 _12202_ ( .A1(_04775_ ), .A2(_04792_ ), .A3(_04794_ ), .A4(_04797_ ), .ZN(_04798_ ) );
NAND2_X1 _12203_ ( .A1(_04535_ ), .A2(fanout_net_16 ), .ZN(_04799_ ) );
NAND3_X1 _12204_ ( .A1(_04519_ ), .A2(_04524_ ), .A3(_04495_ ), .ZN(_04800_ ) );
NAND2_X1 _12205_ ( .A1(_04799_ ), .A2(_04800_ ), .ZN(_04801_ ) );
AOI21_X1 _12206_ ( .A(fanout_net_17 ), .B1(_04571_ ), .B2(_04574_ ), .ZN(_04802_ ) );
AOI21_X1 _12207_ ( .A(_04494_ ), .B1(_04511_ ), .B2(_04514_ ), .ZN(_04803_ ) );
NOR2_X1 _12208_ ( .A1(_04802_ ), .A2(_04803_ ), .ZN(_04804_ ) );
MUX2_X1 _12209_ ( .A(_04801_ ), .B(_04804_ ), .S(_04754_ ), .Z(_04805_ ) );
AOI21_X1 _12210_ ( .A(_03079_ ), .B1(_04805_ ), .B2(_04757_ ), .ZN(_04806_ ) );
AOI211_X1 _12211_ ( .A(_04460_ ), .B(_04770_ ), .C1(_04798_ ), .C2(_04806_ ), .ZN(_00308_ ) );
AND4_X1 _12212_ ( .A1(_03324_ ), .A2(_04486_ ), .A3(_04487_ ), .A4(fanout_net_19 ), .ZN(_04807_ ) );
NOR2_X1 _12213_ ( .A1(_04643_ ), .A2(fanout_net_17 ), .ZN(_04808_ ) );
NAND3_X1 _12214_ ( .A1(_04808_ ), .A2(_04630_ ), .A3(_04505_ ), .ZN(_04809_ ) );
NAND2_X1 _12215_ ( .A1(_03113_ ), .A2(_03482_ ), .ZN(_04810_ ) );
AOI21_X1 _12216_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [18] ), .B2(\u_exu.alu_p2 [18] ), .ZN(_04811_ ) );
OAI211_X1 _12217_ ( .A(_03401_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [18] ), .C2(\u_exu.alu_p2 [18] ), .ZN(_04812_ ) );
OAI211_X1 _12218_ ( .A(_04809_ ), .B(_04810_ ), .C1(_04811_ ), .C2(_04812_ ), .ZN(_04813_ ) );
OAI211_X1 _12219_ ( .A(_03452_ ), .B(_03470_ ), .C1(\u_exu.alu_p2 [0] ), .C2(_03299_ ), .ZN(_04814_ ) );
NAND3_X1 _12220_ ( .A1(_03469_ ), .A2(fanout_net_15 ), .A3(_03472_ ), .ZN(_04815_ ) );
AND2_X1 _12221_ ( .A1(_04814_ ), .A2(_04815_ ), .ZN(_04816_ ) );
OR3_X1 _12222_ ( .A1(_03448_ ), .A2(_03449_ ), .A3(_03096_ ), .ZN(_04817_ ) );
OR3_X1 _12223_ ( .A1(_03440_ ), .A2(_03441_ ), .A3(fanout_net_15 ), .ZN(_04818_ ) );
AND2_X1 _12224_ ( .A1(_04817_ ), .A2(_04818_ ), .ZN(_04819_ ) );
MUX2_X1 _12225_ ( .A(_04816_ ), .B(_04819_ ), .S(_03101_ ), .Z(_04820_ ) );
AND2_X1 _12226_ ( .A1(_04820_ ), .A2(_04493_ ), .ZN(_04821_ ) );
OR3_X1 _12227_ ( .A1(_03460_ ), .A2(_03100_ ), .A3(fanout_net_15 ), .ZN(_04822_ ) );
NOR2_X1 _12228_ ( .A1(_03463_ ), .A2(_03465_ ), .ZN(_04823_ ) );
MUX2_X1 _12229_ ( .A(_04823_ ), .B(_03459_ ), .S(fanout_net_15 ), .Z(_04824_ ) );
OAI21_X1 _12230_ ( .A(_04822_ ), .B1(_04824_ ), .B2(fanout_net_17 ), .ZN(_04825_ ) );
AND2_X1 _12231_ ( .A1(_04825_ ), .A2(fanout_net_18 ), .ZN(_04826_ ) );
NOR2_X1 _12232_ ( .A1(_04821_ ), .A2(_04826_ ), .ZN(_04827_ ) );
AOI21_X1 _12233_ ( .A(_04825_ ), .B1(fanout_net_15 ), .B2(_04678_ ), .ZN(_04828_ ) );
NOR2_X1 _12234_ ( .A1(_04828_ ), .A2(_04507_ ), .ZN(_04829_ ) );
NOR2_X1 _12235_ ( .A1(_04829_ ), .A2(_04821_ ), .ZN(_04830_ ) );
OAI221_X1 _12236_ ( .A(_04677_ ), .B1(_04827_ ), .B2(_04732_ ), .C1(_04830_ ), .C2(_04684_ ), .ZN(_04831_ ) );
NOR4_X1 _12237_ ( .A1(_04772_ ), .A2(_04723_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03490_ ), .ZN(_04832_ ) );
NAND3_X1 _12238_ ( .A1(_04771_ ), .A2(_03332_ ), .A3(_03331_ ), .ZN(_04833_ ) );
AOI221_X4 _12239_ ( .A(_04813_ ), .B1(_04737_ ), .B2(_04831_ ), .C1(_04832_ ), .C2(_04833_ ), .ZN(_04834_ ) );
NAND3_X1 _12240_ ( .A1(_04631_ ), .A2(_04632_ ), .A3(_04516_ ), .ZN(_04835_ ) );
NAND3_X1 _12241_ ( .A1(_04638_ ), .A2(_04639_ ), .A3(fanout_net_17 ), .ZN(_04836_ ) );
NAND3_X1 _12242_ ( .A1(_04835_ ), .A2(_04836_ ), .A3(fanout_net_18 ), .ZN(_04837_ ) );
NAND2_X1 _12243_ ( .A1(_04634_ ), .A2(_04635_ ), .ZN(_04838_ ) );
NAND2_X1 _12244_ ( .A1(_04838_ ), .A2(fanout_net_17 ), .ZN(_04839_ ) );
NAND3_X1 _12245_ ( .A1(_04623_ ), .A2(_04624_ ), .A3(_04538_ ), .ZN(_04840_ ) );
NAND3_X1 _12246_ ( .A1(_04839_ ), .A2(_04840_ ), .A3(_04754_ ), .ZN(_04841_ ) );
NAND3_X1 _12247_ ( .A1(_04837_ ), .A2(_04841_ ), .A3(_04757_ ), .ZN(_04842_ ) );
AND2_X1 _12248_ ( .A1(_04842_ ), .A2(_04653_ ), .ZN(_04843_ ) );
AOI211_X1 _12249_ ( .A(_04460_ ), .B(_04807_ ), .C1(_04834_ ), .C2(_04843_ ), .ZN(_00309_ ) );
NOR2_X1 _12250_ ( .A1(_03312_ ), .A2(\u_exu.alu_p1 [16] ), .ZN(_04844_ ) );
NOR3_X1 _12251_ ( .A1(_03291_ ), .A2(_03328_ ), .A3(_04844_ ), .ZN(_04845_ ) );
OR3_X1 _12252_ ( .A1(_04845_ ), .A2(_03317_ ), .A3(_03328_ ), .ZN(_04846_ ) );
OAI21_X1 _12253_ ( .A(_03317_ ), .B1(_04845_ ), .B2(_03328_ ), .ZN(_04847_ ) );
AND3_X1 _12254_ ( .A1(_04846_ ), .A2(_04549_ ), .A3(_04847_ ), .ZN(_04848_ ) );
MUX2_X1 _12255_ ( .A(_04674_ ), .B(_04669_ ), .S(_03101_ ), .Z(_04849_ ) );
NOR2_X1 _12256_ ( .A1(_04849_ ), .A2(_04629_ ), .ZN(_04850_ ) );
AOI21_X1 _12257_ ( .A(_03101_ ), .B1(_04663_ ), .B2(_04664_ ), .ZN(_04851_ ) );
OAI21_X1 _12258_ ( .A(_04527_ ), .B1(_04569_ ), .B2(_04573_ ), .ZN(_04852_ ) );
OAI21_X1 _12259_ ( .A(fanout_net_15 ), .B1(_04572_ ), .B2(_04578_ ), .ZN(_04853_ ) );
AND3_X1 _12260_ ( .A1(_04852_ ), .A2(_04853_ ), .A3(_03101_ ), .ZN(_04854_ ) );
NOR3_X1 _12261_ ( .A1(_04851_ ), .A2(_04854_ ), .A3(fanout_net_18 ), .ZN(_04855_ ) );
OAI21_X1 _12262_ ( .A(_04608_ ), .B1(_04850_ ), .B2(_04855_ ), .ZN(_04856_ ) );
AND2_X1 _12263_ ( .A1(_04856_ ), .A2(_04677_ ), .ZN(_04857_ ) );
OR2_X1 _12264_ ( .A1(_04680_ ), .A2(_04494_ ), .ZN(_04858_ ) );
OAI21_X1 _12265_ ( .A(_04858_ ), .B1(fanout_net_17 ), .B2(_04669_ ), .ZN(_04859_ ) );
AND2_X1 _12266_ ( .A1(_04859_ ), .A2(fanout_net_18 ), .ZN(_04860_ ) );
OAI21_X1 _12267_ ( .A(_04599_ ), .B1(_04860_ ), .B2(_04855_ ), .ZN(_04861_ ) );
AOI21_X1 _12268_ ( .A(_03437_ ), .B1(_04857_ ), .B2(_04861_ ), .ZN(_04862_ ) );
NAND2_X1 _12269_ ( .A1(_04694_ ), .A2(_04516_ ), .ZN(_04863_ ) );
NAND2_X1 _12270_ ( .A1(_04704_ ), .A2(fanout_net_17 ), .ZN(_04864_ ) );
CLKBUF_X2 _12271_ ( .A(_04493_ ), .Z(_04865_ ) );
AND3_X1 _12272_ ( .A1(_04863_ ), .A2(_04864_ ), .A3(_04865_ ), .ZN(_04866_ ) );
AOI21_X1 _12273_ ( .A(fanout_net_17 ), .B1(_04697_ ), .B2(_04698_ ), .ZN(_04867_ ) );
AOI21_X1 _12274_ ( .A(_04537_ ), .B1(_04711_ ), .B2(_04712_ ), .ZN(_04868_ ) );
CLKBUF_X2 _12275_ ( .A(_04493_ ), .Z(_04869_ ) );
NOR3_X1 _12276_ ( .A1(_04867_ ), .A2(_04868_ ), .A3(_04869_ ), .ZN(_04870_ ) );
NOR3_X1 _12277_ ( .A1(_04866_ ), .A2(_04870_ ), .A3(_04589_ ), .ZN(_04871_ ) );
NOR3_X1 _12278_ ( .A1(_04709_ ), .A2(fanout_net_17 ), .A3(fanout_net_15 ), .ZN(_04872_ ) );
NAND3_X1 _12279_ ( .A1(_04872_ ), .A2(_04630_ ), .A3(_04505_ ), .ZN(_04873_ ) );
NAND2_X1 _12280_ ( .A1(_03112_ ), .A2(_03482_ ), .ZN(_04874_ ) );
AOI21_X1 _12281_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p2 [17] ), .B2(\u_exu.alu_p1 [17] ), .ZN(_04875_ ) );
OAI211_X1 _12282_ ( .A(_03401_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p2 [17] ), .C2(\u_exu.alu_p1 [17] ), .ZN(_04876_ ) );
OAI211_X1 _12283_ ( .A(_04873_ ), .B(_04874_ ), .C1(_04875_ ), .C2(_04876_ ), .ZN(_04877_ ) );
OR4_X1 _12284_ ( .A1(_04848_ ), .A2(_04862_ ), .A3(_04871_ ), .A4(_04877_ ), .ZN(_04878_ ) );
BUF_X4 _12285_ ( .A(_04653_ ), .Z(_04879_ ) );
MUX2_X1 _12286_ ( .A(\u_exu.alu_p1 [17] ), .B(_04878_ ), .S(_04879_ ), .Z(_04880_ ) );
AND2_X1 _12287_ ( .A1(_04880_ ), .A2(_04593_ ), .ZN(_00310_ ) );
NOR4_X1 _12288_ ( .A1(_04845_ ), .A2(_04723_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03490_ ), .ZN(_04881_ ) );
OAI21_X1 _12289_ ( .A(_04881_ ), .B1(_03292_ ), .B2(_03314_ ), .ZN(_04882_ ) );
NOR4_X1 _12290_ ( .A1(_03153_ ), .A2(_04723_ ), .A3(_04486_ ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_04883_ ) );
OAI21_X1 _12291_ ( .A(_04883_ ), .B1(fanout_net_11 ), .B2(_03152_ ), .ZN(_04884_ ) );
INV_X1 _12292_ ( .A(_04767_ ), .ZN(_04885_ ) );
OR3_X1 _12293_ ( .A1(_04885_ ), .A2(_03153_ ), .A3(_03152_ ), .ZN(_04886_ ) );
NOR2_X1 _12294_ ( .A1(_03476_ ), .A2(\u_exu.alu_p2 [4] ), .ZN(_04887_ ) );
OAI21_X1 _12295_ ( .A(_04737_ ), .B1(_04887_ ), .B2(_04606_ ), .ZN(_04888_ ) );
NAND2_X1 _12296_ ( .A1(_04741_ ), .A2(_04538_ ), .ZN(_04889_ ) );
NAND2_X1 _12297_ ( .A1(_04761_ ), .A2(fanout_net_17 ), .ZN(_04890_ ) );
NAND3_X1 _12298_ ( .A1(_04889_ ), .A2(_04890_ ), .A3(fanout_net_18 ), .ZN(_04891_ ) );
NAND2_X1 _12299_ ( .A1(_04749_ ), .A2(_04538_ ), .ZN(_04892_ ) );
NAND3_X1 _12300_ ( .A1(_04743_ ), .A2(_04744_ ), .A3(fanout_net_17 ), .ZN(_04893_ ) );
NAND3_X1 _12301_ ( .A1(_04892_ ), .A2(_04893_ ), .A3(_04754_ ), .ZN(_04894_ ) );
NAND3_X1 _12302_ ( .A1(_04891_ ), .A2(_04894_ ), .A3(_04757_ ), .ZN(_04895_ ) );
AND3_X1 _12303_ ( .A1(_03095_ ), .A2(_04537_ ), .A3(_04491_ ), .ZN(_04896_ ) );
NAND3_X1 _12304_ ( .A1(_04506_ ), .A2(_04754_ ), .A3(_04896_ ), .ZN(_04897_ ) );
AND3_X1 _12305_ ( .A1(_04888_ ), .A2(_04895_ ), .A3(_04897_ ), .ZN(_04898_ ) );
NAND4_X1 _12306_ ( .A1(_04882_ ), .A2(_04884_ ), .A3(_04886_ ), .A4(_04898_ ), .ZN(_04899_ ) );
BUF_X4 _12307_ ( .A(_04653_ ), .Z(_04900_ ) );
MUX2_X1 _12308_ ( .A(\u_exu.alu_p1 [16] ), .B(_04899_ ), .S(_04900_ ), .Z(_04901_ ) );
AND2_X1 _12309_ ( .A1(_04901_ ), .A2(_04593_ ), .ZN(_00311_ ) );
NOR4_X1 _12310_ ( .A1(_04724_ ), .A2(\u_exu.alu_p1 [15] ), .A3(\u_exu.alu_ctrl [5] ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_04902_ ) );
INV_X1 _12311_ ( .A(_03225_ ), .ZN(_04903_ ) );
INV_X1 _12312_ ( .A(_03219_ ), .ZN(_04904_ ) );
OAI21_X1 _12313_ ( .A(_03243_ ), .B1(_03282_ ), .B2(_03289_ ), .ZN(_04905_ ) );
AOI21_X1 _12314_ ( .A(_04904_ ), .B1(_04905_ ), .B2(_03215_ ), .ZN(_04906_ ) );
XNOR2_X1 _12315_ ( .A(_03220_ ), .B(_03170_ ), .ZN(_04907_ ) );
OAI22_X1 _12316_ ( .A1(_04906_ ), .A2(_03234_ ), .B1(\u_exu.alu_p1 [13] ), .B2(_04907_ ), .ZN(_04908_ ) );
AOI21_X1 _12317_ ( .A(_04903_ ), .B1(_04908_ ), .B2(_03233_ ), .ZN(_04909_ ) );
OR3_X1 _12318_ ( .A1(_04909_ ), .A2(_03187_ ), .A3(_03190_ ), .ZN(_04910_ ) );
OAI21_X1 _12319_ ( .A(_03187_ ), .B1(_04909_ ), .B2(_03190_ ), .ZN(_04911_ ) );
NAND3_X1 _12320_ ( .A1(_04910_ ), .A2(_04550_ ), .A3(_04911_ ), .ZN(_04912_ ) );
NAND2_X1 _12321_ ( .A1(_03136_ ), .A2(_04767_ ), .ZN(_04913_ ) );
AOI21_X1 _12322_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [15] ), .B2(\u_exu.alu_p2 [15] ), .ZN(_04914_ ) );
OAI211_X1 _12323_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [15] ), .C2(\u_exu.alu_p2 [15] ), .ZN(_04915_ ) );
OAI211_X1 _12324_ ( .A(_04913_ ), .B(_04653_ ), .C1(_04914_ ), .C2(_04915_ ), .ZN(_04916_ ) );
BUF_X4 _12325_ ( .A(_04618_ ), .Z(_04917_ ) );
NAND3_X1 _12326_ ( .A1(_04783_ ), .A2(_04784_ ), .A3(_04495_ ), .ZN(_04918_ ) );
OAI21_X1 _12327_ ( .A(_04918_ ), .B1(_04777_ ), .B2(_04537_ ), .ZN(_04919_ ) );
AND2_X1 _12328_ ( .A1(_04919_ ), .A2(fanout_net_18 ), .ZN(_04920_ ) );
OR3_X1 _12329_ ( .A1(_04569_ ), .A2(_04527_ ), .A3(_04573_ ), .ZN(_04921_ ) );
OR3_X1 _12330_ ( .A1(_04509_ ), .A2(fanout_net_15 ), .A3(_04570_ ), .ZN(_04922_ ) );
NAND2_X1 _12331_ ( .A1(_04921_ ), .A2(_04922_ ), .ZN(_04923_ ) );
NAND2_X1 _12332_ ( .A1(_04923_ ), .A2(_04537_ ), .ZN(_04924_ ) );
NAND2_X1 _12333_ ( .A1(_04780_ ), .A2(_04781_ ), .ZN(_04925_ ) );
NAND2_X1 _12334_ ( .A1(_04925_ ), .A2(fanout_net_17 ), .ZN(_04926_ ) );
AND3_X1 _12335_ ( .A1(_04924_ ), .A2(_04926_ ), .A3(_04508_ ), .ZN(_04927_ ) );
OAI21_X1 _12336_ ( .A(_04917_ ), .B1(_04920_ ), .B2(_04927_ ), .ZN(_04928_ ) );
NAND3_X1 _12337_ ( .A1(_04489_ ), .A2(_04495_ ), .A3(_04491_ ), .ZN(_04929_ ) );
NOR2_X1 _12338_ ( .A1(_03098_ ), .A2(\u_exu.alu_ctrl [1] ), .ZN(_04930_ ) );
INV_X1 _12339_ ( .A(_04930_ ), .ZN(_04931_ ) );
NOR3_X1 _12340_ ( .A1(_04929_ ), .A2(fanout_net_18 ), .A3(_04931_ ), .ZN(_04932_ ) );
NOR2_X1 _12341_ ( .A1(_04932_ ), .A2(_04606_ ), .ZN(_04933_ ) );
AOI21_X1 _12342_ ( .A(_03437_ ), .B1(_04928_ ), .B2(_04933_ ), .ZN(_04934_ ) );
AOI211_X1 _12343_ ( .A(_04916_ ), .B(_04934_ ), .C1(_04546_ ), .C2(_04757_ ), .ZN(_04935_ ) );
AOI211_X1 _12344_ ( .A(_04460_ ), .B(_04902_ ), .C1(_04912_ ), .C2(_04935_ ), .ZN(_00312_ ) );
AND4_X1 _12345_ ( .A1(_03224_ ), .A2(_04486_ ), .A3(_04487_ ), .A4(fanout_net_19 ), .ZN(_04936_ ) );
NOR4_X1 _12346_ ( .A1(_04909_ ), .A2(_04724_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_04487_ ), .ZN(_04937_ ) );
NAND3_X1 _12347_ ( .A1(_04908_ ), .A2(_04903_ ), .A3(_03233_ ), .ZN(_04938_ ) );
NAND2_X1 _12348_ ( .A1(_04937_ ), .A2(_04938_ ), .ZN(_04939_ ) );
INV_X1 _12349_ ( .A(_04605_ ), .ZN(_04940_ ) );
OR3_X1 _12350_ ( .A1(_04602_ ), .A2(_04603_ ), .A3(_04940_ ), .ZN(_04941_ ) );
OAI211_X1 _12351_ ( .A(_04941_ ), .B(_04737_ ), .C1(_04607_ ), .C2(_04931_ ), .ZN(_04942_ ) );
NOR2_X1 _12352_ ( .A1(_04824_ ), .A2(_03101_ ), .ZN(_04943_ ) );
AOI21_X1 _12353_ ( .A(_04943_ ), .B1(_03102_ ), .B2(_04816_ ), .ZN(_04944_ ) );
NOR2_X1 _12354_ ( .A1(_04944_ ), .A2(_04754_ ), .ZN(_04945_ ) );
AOI21_X1 _12355_ ( .A(_03102_ ), .B1(_04817_ ), .B2(_04818_ ), .ZN(_04946_ ) );
OR3_X1 _12356_ ( .A1(_03443_ ), .A2(_03444_ ), .A3(_04490_ ), .ZN(_04947_ ) );
OR3_X1 _12357_ ( .A1(_03426_ ), .A2(_03427_ ), .A3(fanout_net_15 ), .ZN(_04948_ ) );
AOI21_X1 _12358_ ( .A(fanout_net_17 ), .B1(_04947_ ), .B2(_04948_ ), .ZN(_04949_ ) );
NOR2_X1 _12359_ ( .A1(_04946_ ), .A2(_04949_ ), .ZN(_04950_ ) );
AOI21_X1 _12360_ ( .A(_04945_ ), .B1(_04754_ ), .B2(_04950_ ), .ZN(_04951_ ) );
AOI21_X1 _12361_ ( .A(_04942_ ), .B1(_04951_ ), .B2(_04917_ ), .ZN(_04952_ ) );
AND3_X1 _12362_ ( .A1(_04637_ ), .A2(_04644_ ), .A3(_04757_ ), .ZN(_04953_ ) );
NAND2_X1 _12363_ ( .A1(_03118_ ), .A2(_04767_ ), .ZN(_04954_ ) );
AOI21_X1 _12364_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [14] ), .B2(\u_exu.alu_p2 [14] ), .ZN(_04955_ ) );
OAI211_X1 _12365_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [14] ), .C2(\u_exu.alu_p2 [14] ), .ZN(_04956_ ) );
OAI211_X1 _12366_ ( .A(_04954_ ), .B(_04653_ ), .C1(_04955_ ), .C2(_04956_ ), .ZN(_04957_ ) );
NOR3_X1 _12367_ ( .A1(_04952_ ), .A2(_04953_ ), .A3(_04957_ ), .ZN(_04958_ ) );
AOI211_X1 _12368_ ( .A(_04460_ ), .B(_04936_ ), .C1(_04939_ ), .C2(_04958_ ), .ZN(_00313_ ) );
OR3_X1 _12369_ ( .A1(_04906_ ), .A2(_03234_ ), .A3(_03222_ ), .ZN(_04959_ ) );
OAI21_X1 _12370_ ( .A(_03222_ ), .B1(_04906_ ), .B2(_03234_ ), .ZN(_04960_ ) );
NAND3_X1 _12371_ ( .A1(_04959_ ), .A2(_04549_ ), .A3(_04960_ ), .ZN(_04961_ ) );
OR2_X1 _12372_ ( .A1(_04714_ ), .A2(_04493_ ), .ZN(_04962_ ) );
NAND3_X1 _12373_ ( .A1(_04700_ ), .A2(_04705_ ), .A3(_04629_ ), .ZN(_04963_ ) );
AND3_X1 _12374_ ( .A1(_04962_ ), .A2(_04588_ ), .A3(_04963_ ), .ZN(_04964_ ) );
NAND2_X1 _12375_ ( .A1(_04670_ ), .A2(fanout_net_18 ), .ZN(_04965_ ) );
OR3_X1 _12376_ ( .A1(_04509_ ), .A2(_03470_ ), .A3(_04570_ ), .ZN(_04966_ ) );
OR3_X1 _12377_ ( .A1(_04702_ ), .A2(_04510_ ), .A3(fanout_net_15 ), .ZN(_04967_ ) );
AOI21_X1 _12378_ ( .A(fanout_net_17 ), .B1(_04966_ ), .B2(_04967_ ), .ZN(_04968_ ) );
AND3_X1 _12379_ ( .A1(_04852_ ), .A2(_04853_ ), .A3(fanout_net_17 ), .ZN(_04969_ ) );
OR2_X1 _12380_ ( .A1(_04968_ ), .A2(_04969_ ), .ZN(_04970_ ) );
OAI211_X1 _12381_ ( .A(_04965_ ), .B(_04917_ ), .C1(fanout_net_18 ), .C2(_04970_ ), .ZN(_04971_ ) );
NOR2_X1 _12382_ ( .A1(_04603_ ), .A2(_04497_ ), .ZN(_04972_ ) );
INV_X1 _12383_ ( .A(_04972_ ), .ZN(_04973_ ) );
AOI21_X1 _12384_ ( .A(_04973_ ), .B1(_04681_ ), .B2(_04629_ ), .ZN(_04974_ ) );
NOR2_X1 _12385_ ( .A1(_04674_ ), .A2(fanout_net_17 ), .ZN(_04975_ ) );
NAND3_X1 _12386_ ( .A1(_04975_ ), .A2(_04629_ ), .A3(_04686_ ), .ZN(_04976_ ) );
AND2_X1 _12387_ ( .A1(_04686_ ), .A2(_04931_ ), .ZN(_04977_ ) );
INV_X1 _12388_ ( .A(_04977_ ), .ZN(_04978_ ) );
AOI22_X1 _12389_ ( .A1(_04974_ ), .A2(\u_exu.alu_p2 [4] ), .B1(_04976_ ), .B2(_04978_ ), .ZN(_04979_ ) );
AOI221_X4 _12390_ ( .A(_04964_ ), .B1(_03119_ ), .B2(_03482_ ), .C1(_04971_ ), .C2(_04979_ ), .ZN(_04980_ ) );
AOI21_X1 _12391_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [13] ), .B2(\u_exu.alu_p2 [13] ), .ZN(_04981_ ) );
BUF_X4 _12392_ ( .A(_04649_ ), .Z(_04982_ ) );
OAI211_X1 _12393_ ( .A(_04982_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [13] ), .C2(\u_exu.alu_p2 [13] ), .ZN(_04983_ ) );
OAI211_X1 _12394_ ( .A(_04961_ ), .B(_04980_ ), .C1(_04981_ ), .C2(_04983_ ), .ZN(_04984_ ) );
MUX2_X1 _12395_ ( .A(\u_exu.alu_p1 [13] ), .B(_04984_ ), .S(_04879_ ), .Z(_04985_ ) );
AND2_X1 _12396_ ( .A1(_04985_ ), .A2(_04593_ ), .ZN(_00314_ ) );
NOR4_X1 _12397_ ( .A1(_04906_ ), .A2(_04724_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03490_ ), .ZN(_04986_ ) );
NAND3_X1 _12398_ ( .A1(_04905_ ), .A2(_04904_ ), .A3(_03215_ ), .ZN(_04987_ ) );
NAND2_X1 _12399_ ( .A1(_04986_ ), .A2(_04987_ ), .ZN(_04988_ ) );
AND2_X1 _12400_ ( .A1(_04762_ ), .A2(\u_exu.alu_p2 [3] ), .ZN(_04989_ ) );
AOI21_X1 _12401_ ( .A(\u_exu.alu_p2 [3] ), .B1(_04742_ ), .B2(_04745_ ), .ZN(_04990_ ) );
NOR2_X1 _12402_ ( .A1(_04989_ ), .A2(_04990_ ), .ZN(_04991_ ) );
NOR2_X1 _12403_ ( .A1(_04991_ ), .A2(_04589_ ), .ZN(_04992_ ) );
NOR2_X1 _12404_ ( .A1(_03461_ ), .A2(fanout_net_17 ), .ZN(_04993_ ) );
NAND3_X1 _12405_ ( .A1(_04993_ ), .A2(_04630_ ), .A3(_04686_ ), .ZN(_04994_ ) );
NAND2_X1 _12406_ ( .A1(_04994_ ), .A2(_04978_ ), .ZN(_04995_ ) );
OR2_X1 _12407_ ( .A1(_04728_ ), .A2(_04507_ ), .ZN(_04996_ ) );
NAND3_X1 _12408_ ( .A1(_03428_ ), .A2(_03431_ ), .A3(_04494_ ), .ZN(_04997_ ) );
OAI21_X1 _12409_ ( .A(_04997_ ), .B1(_03446_ ), .B2(_03102_ ), .ZN(_04998_ ) );
AOI21_X1 _12410_ ( .A(\u_exu.alu_p2 [4] ), .B1(_04998_ ), .B2(_04865_ ), .ZN(_04999_ ) );
AOI21_X1 _12411_ ( .A(_04973_ ), .B1(_04733_ ), .B2(_04865_ ), .ZN(_05000_ ) );
AOI22_X1 _12412_ ( .A1(_04996_ ), .A2(_04999_ ), .B1(\u_exu.alu_p2 [4] ), .B2(_05000_ ), .ZN(_05001_ ) );
AOI221_X4 _12413_ ( .A(_04992_ ), .B1(_03134_ ), .B2(_04646_ ), .C1(_04995_ ), .C2(_05001_ ), .ZN(_05002_ ) );
AOI21_X1 _12414_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [12] ), .B2(\u_exu.alu_p2 [12] ), .ZN(_05003_ ) );
OAI211_X1 _12415_ ( .A(_04982_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [12] ), .C2(\u_exu.alu_p2 [12] ), .ZN(_05004_ ) );
OAI211_X1 _12416_ ( .A(_04988_ ), .B(_05002_ ), .C1(_05003_ ), .C2(_05004_ ), .ZN(_05005_ ) );
MUX2_X1 _12417_ ( .A(\u_exu.alu_p1 [12] ), .B(_05005_ ), .S(_04900_ ), .Z(_05006_ ) );
AND2_X1 _12418_ ( .A1(_05006_ ), .A2(_04593_ ), .ZN(_00315_ ) );
AOI21_X1 _12419_ ( .A(_03184_ ), .B1(_03369_ ), .B2(_03381_ ), .ZN(_05007_ ) );
OR3_X4 _12420_ ( .A1(_05007_ ), .A2(_03178_ ), .A3(_03383_ ), .ZN(_05008_ ) );
OAI21_X1 _12421_ ( .A(_03178_ ), .B1(_05007_ ), .B2(_03383_ ), .ZN(_05009_ ) );
AND3_X2 _12422_ ( .A1(_05008_ ), .A2(_04549_ ), .A3(_05009_ ), .ZN(_05010_ ) );
OAI211_X1 _12423_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [29] ), .C2(\u_exu.alu_p2 [29] ), .ZN(_05011_ ) );
AOI21_X1 _12424_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [29] ), .B2(\u_exu.alu_p2 [29] ), .ZN(_05012_ ) );
NOR2_X1 _12425_ ( .A1(_05011_ ), .A2(_05012_ ), .ZN(_05013_ ) );
AND2_X1 _12426_ ( .A1(_03123_ ), .A2(_04646_ ), .ZN(_05014_ ) );
NAND3_X1 _12427_ ( .A1(_04962_ ), .A2(_04506_ ), .A3(_04963_ ), .ZN(_05015_ ) );
NAND3_X1 _12428_ ( .A1(_04691_ ), .A2(_04695_ ), .A3(\u_exu.alu_p2 [3] ), .ZN(_05016_ ) );
OR3_X1 _12429_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(fanout_net_15 ), .ZN(_05017_ ) );
OAI211_X1 _12430_ ( .A(_04559_ ), .B(fanout_net_15 ), .C1(\u_exu.alu_p2 [0] ), .C2(_03355_ ), .ZN(_05018_ ) );
NAND3_X1 _12431_ ( .A1(_05017_ ), .A2(_05018_ ), .A3(_04516_ ), .ZN(_05019_ ) );
NAND3_X1 _12432_ ( .A1(_04582_ ), .A2(fanout_net_15 ), .A3(_04584_ ), .ZN(_05020_ ) );
NAND3_X1 _12433_ ( .A1(_04562_ ), .A2(_04491_ ), .A3(_04564_ ), .ZN(_05021_ ) );
NAND2_X1 _12434_ ( .A1(_05020_ ), .A2(_05021_ ), .ZN(_05022_ ) );
OAI211_X1 _12435_ ( .A(_05019_ ), .B(_04869_ ), .C1(_04538_ ), .C2(_05022_ ), .ZN(_05023_ ) );
NAND3_X1 _12436_ ( .A1(_05016_ ), .A2(_04756_ ), .A3(_05023_ ), .ZN(_05024_ ) );
MUX2_X1 _12437_ ( .A(_03395_ ), .B(_04974_ ), .S(_04618_ ), .Z(_05025_ ) );
AND2_X1 _12438_ ( .A1(_04975_ ), .A2(_04865_ ), .ZN(_05026_ ) );
OAI21_X1 _12439_ ( .A(_04977_ ), .B1(_05026_ ), .B2(\u_exu.alu_ctrl [1] ), .ZN(_05027_ ) );
OAI211_X1 _12440_ ( .A(_05015_ ), .B(_05024_ ), .C1(_05025_ ), .C2(_05027_ ), .ZN(_05028_ ) );
OR4_X4 _12441_ ( .A1(_05010_ ), .A2(_05013_ ), .A3(_05014_ ), .A4(_05028_ ), .ZN(_05029_ ) );
MUX2_X2 _12442_ ( .A(\u_exu.alu_p1 [29] ), .B(_05029_ ), .S(_04900_ ), .Z(_05030_ ) );
AND2_X1 _12443_ ( .A1(_05030_ ), .A2(_04593_ ), .ZN(_00316_ ) );
NOR4_X1 _12444_ ( .A1(_04724_ ), .A2(\u_exu.alu_p1 [11] ), .A3(\u_exu.alu_ctrl [5] ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_05031_ ) );
OAI21_X1 _12445_ ( .A(_03242_ ), .B1(_03282_ ), .B2(_03289_ ), .ZN(_05032_ ) );
AOI21_X1 _12446_ ( .A(_03205_ ), .B1(_05032_ ), .B2(_03200_ ), .ZN(_05033_ ) );
OR3_X1 _12447_ ( .A1(_05033_ ), .A2(_03212_ ), .A3(_03213_ ), .ZN(_05034_ ) );
OAI21_X1 _12448_ ( .A(_03212_ ), .B1(_05033_ ), .B2(_03213_ ), .ZN(_05035_ ) );
NAND3_X1 _12449_ ( .A1(_05034_ ), .A2(_04550_ ), .A3(_05035_ ), .ZN(_05036_ ) );
NAND3_X1 _12450_ ( .A1(_04799_ ), .A2(_04800_ ), .A3(_04507_ ), .ZN(_05037_ ) );
OAI21_X1 _12451_ ( .A(\u_exu.alu_p2 [3] ), .B1(_04544_ ), .B2(fanout_net_17 ), .ZN(_05038_ ) );
NAND3_X1 _12452_ ( .A1(_05037_ ), .A2(_05038_ ), .A3(_04757_ ), .ZN(_05039_ ) );
AOI21_X1 _12453_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [11] ), .B2(\u_exu.alu_p2 [11] ), .ZN(_05040_ ) );
OAI211_X1 _12454_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [11] ), .C2(\u_exu.alu_p2 [11] ), .ZN(_05041_ ) );
AOI21_X1 _12455_ ( .A(\u_exu.alu_p2 [3] ), .B1(_04789_ ), .B2(_04679_ ), .ZN(_05042_ ) );
NOR2_X1 _12456_ ( .A1(_05042_ ), .A2(_04973_ ), .ZN(_05043_ ) );
NAND2_X1 _12457_ ( .A1(_04923_ ), .A2(fanout_net_17 ), .ZN(_05044_ ) );
OAI21_X1 _12458_ ( .A(_04528_ ), .B1(_04520_ ), .B2(_04512_ ), .ZN(_05045_ ) );
OAI21_X1 _12459_ ( .A(\u_exu.alu_p2 [1] ), .B1(_04702_ ), .B2(_04510_ ), .ZN(_05046_ ) );
NAND3_X1 _12460_ ( .A1(_05045_ ), .A2(_03102_ ), .A3(_05046_ ), .ZN(_05047_ ) );
NAND2_X1 _12461_ ( .A1(_05044_ ), .A2(_05047_ ), .ZN(_05048_ ) );
OR2_X1 _12462_ ( .A1(_04782_ ), .A2(_04785_ ), .ZN(_05049_ ) );
MUX2_X1 _12463_ ( .A(_05048_ ), .B(_05049_ ), .S(\u_exu.alu_p2 [3] ), .Z(_05050_ ) );
MUX2_X1 _12464_ ( .A(_05043_ ), .B(_05050_ ), .S(_04917_ ), .Z(_05051_ ) );
NAND3_X1 _12465_ ( .A1(_04778_ ), .A2(_04508_ ), .A3(_04686_ ), .ZN(_05052_ ) );
AND2_X1 _12466_ ( .A1(_05052_ ), .A2(_04978_ ), .ZN(_05053_ ) );
OAI221_X1 _12467_ ( .A(_05039_ ), .B1(_05040_ ), .B2(_05041_ ), .C1(_05051_ ), .C2(_05053_ ), .ZN(_05054_ ) );
AOI211_X1 _12468_ ( .A(_03079_ ), .B(_05054_ ), .C1(_03116_ ), .C2(_04767_ ), .ZN(_05055_ ) );
AOI211_X1 _12469_ ( .A(_04460_ ), .B(_05031_ ), .C1(_05036_ ), .C2(_05055_ ), .ZN(_00317_ ) );
NOR4_X1 _12470_ ( .A1(_05033_ ), .A2(_04723_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03490_ ), .ZN(_05056_ ) );
NAND3_X1 _12471_ ( .A1(_05032_ ), .A2(_03205_ ), .A3(_03200_ ), .ZN(_05057_ ) );
NAND2_X1 _12472_ ( .A1(_05056_ ), .A2(_05057_ ), .ZN(_05058_ ) );
OAI21_X1 _12473_ ( .A(\u_exu.alu_p2 [3] ), .B1(_04643_ ), .B2(fanout_net_17 ), .ZN(_05059_ ) );
NAND3_X1 _12474_ ( .A1(_04835_ ), .A2(_04836_ ), .A3(_04630_ ), .ZN(_05060_ ) );
AND3_X1 _12475_ ( .A1(_05059_ ), .A2(_05060_ ), .A3(_04756_ ), .ZN(_05061_ ) );
OR3_X1 _12476_ ( .A1(_03429_ ), .A2(_03430_ ), .A3(_04527_ ), .ZN(_05062_ ) );
OR3_X1 _12477_ ( .A1(_03419_ ), .A2(_03420_ ), .A3(\u_exu.alu_p2 [1] ), .ZN(_05063_ ) );
NAND3_X1 _12478_ ( .A1(_05062_ ), .A2(_05063_ ), .A3(_03102_ ), .ZN(_05064_ ) );
NAND3_X1 _12479_ ( .A1(_04947_ ), .A2(_04948_ ), .A3(fanout_net_17 ), .ZN(_05065_ ) );
NAND2_X1 _12480_ ( .A1(_05064_ ), .A2(_05065_ ), .ZN(_05066_ ) );
MUX2_X1 _12481_ ( .A(_05066_ ), .B(_04820_ ), .S(\u_exu.alu_p2 [3] ), .Z(_05067_ ) );
AND3_X1 _12482_ ( .A1(_04825_ ), .A2(_04507_ ), .A3(_04686_ ), .ZN(_05068_ ) );
OAI22_X1 _12483_ ( .A1(_05067_ ), .A2(\u_exu.alu_p2 [4] ), .B1(_04977_ ), .B2(_05068_ ), .ZN(_05069_ ) );
NOR2_X1 _12484_ ( .A1(_04828_ ), .A2(\u_exu.alu_p2 [3] ), .ZN(_05070_ ) );
NOR2_X1 _12485_ ( .A1(_05070_ ), .A2(_04973_ ), .ZN(_05071_ ) );
AOI21_X1 _12486_ ( .A(_05069_ ), .B1(\u_exu.alu_p2 [4] ), .B2(_05071_ ), .ZN(_05072_ ) );
AOI211_X1 _12487_ ( .A(_05061_ ), .B(_05072_ ), .C1(_03135_ ), .C2(_04767_ ), .ZN(_05073_ ) );
AOI21_X1 _12488_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [10] ), .B2(\u_exu.alu_p2 [10] ), .ZN(_05074_ ) );
OAI211_X1 _12489_ ( .A(_04982_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [10] ), .C2(\u_exu.alu_p2 [10] ), .ZN(_05075_ ) );
OAI211_X1 _12490_ ( .A(_05058_ ), .B(_05073_ ), .C1(_05074_ ), .C2(_05075_ ), .ZN(_05076_ ) );
MUX2_X1 _12491_ ( .A(\u_exu.alu_p1 [10] ), .B(_05076_ ), .S(_04900_ ), .Z(_05077_ ) );
AND2_X1 _12492_ ( .A1(_05077_ ), .A2(_04593_ ), .ZN(_00318_ ) );
NOR4_X1 _12493_ ( .A1(_04724_ ), .A2(\u_exu.alu_p1 [9] ), .A3(\u_exu.alu_ctrl [5] ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_05078_ ) );
NOR2_X1 _12494_ ( .A1(_03282_ ), .A2(_03289_ ), .ZN(_05079_ ) );
NOR2_X1 _12495_ ( .A1(_03196_ ), .A2(\u_exu.alu_p1 [8] ), .ZN(_05080_ ) );
NOR3_X1 _12496_ ( .A1(_05079_ ), .A2(_03197_ ), .A3(_05080_ ), .ZN(_05081_ ) );
OR3_X1 _12497_ ( .A1(_05081_ ), .A2(_03194_ ), .A3(_03197_ ), .ZN(_05082_ ) );
OAI21_X1 _12498_ ( .A(_03194_ ), .B1(_05081_ ), .B2(_03197_ ), .ZN(_05083_ ) );
NAND3_X1 _12499_ ( .A1(_05082_ ), .A2(_04550_ ), .A3(_05083_ ), .ZN(_05084_ ) );
OAI21_X1 _12500_ ( .A(_04630_ ), .B1(_04867_ ), .B2(_04868_ ), .ZN(_05085_ ) );
NAND3_X1 _12501_ ( .A1(_04710_ ), .A2(\u_exu.alu_p2 [3] ), .A3(_04538_ ), .ZN(_05086_ ) );
AOI21_X1 _12502_ ( .A(_04589_ ), .B1(_05085_ ), .B2(_05086_ ), .ZN(_05087_ ) );
OR3_X1 _12503_ ( .A1(_04851_ ), .A2(_04854_ ), .A3(_03099_ ), .ZN(_05088_ ) );
AOI21_X1 _12504_ ( .A(_03101_ ), .B1(_04966_ ), .B2(_04967_ ), .ZN(_05089_ ) );
OR3_X1 _12505_ ( .A1(_04517_ ), .A2(\u_exu.alu_p2 [1] ), .A3(_04522_ ), .ZN(_05090_ ) );
NAND3_X1 _12506_ ( .A1(_04521_ ), .A2(\u_exu.alu_p2 [1] ), .A3(_04513_ ), .ZN(_05091_ ) );
AOI21_X1 _12507_ ( .A(fanout_net_17 ), .B1(_05090_ ), .B2(_05091_ ), .ZN(_05092_ ) );
NOR2_X1 _12508_ ( .A1(_05089_ ), .A2(_05092_ ), .ZN(_05093_ ) );
AOI21_X1 _12509_ ( .A(\u_exu.alu_p2 [4] ), .B1(_05093_ ), .B2(_04493_ ), .ZN(_05094_ ) );
NOR2_X1 _12510_ ( .A1(_04849_ ), .A2(\u_exu.alu_p2 [3] ), .ZN(_05095_ ) );
INV_X1 _12511_ ( .A(_05095_ ), .ZN(_05096_ ) );
AOI221_X4 _12512_ ( .A(_03437_ ), .B1(_05088_ ), .B2(_05094_ ), .C1(_05096_ ), .C2(_04930_ ), .ZN(_05097_ ) );
AOI21_X1 _12513_ ( .A(_04973_ ), .B1(_04859_ ), .B2(_04630_ ), .ZN(_05098_ ) );
NAND2_X1 _12514_ ( .A1(_05098_ ), .A2(\u_exu.alu_p2 [4] ), .ZN(_05099_ ) );
AOI221_X4 _12515_ ( .A(_05087_ ), .B1(_03139_ ), .B2(_04646_ ), .C1(_05097_ ), .C2(_05099_ ), .ZN(_05100_ ) );
NOR4_X1 _12516_ ( .A1(_03138_ ), .A2(_04724_ ), .A3(_04486_ ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_05101_ ) );
OAI21_X1 _12517_ ( .A(_05101_ ), .B1(fanout_net_11 ), .B2(_03137_ ), .ZN(_05102_ ) );
AND3_X1 _12518_ ( .A1(_05100_ ), .A2(_04879_ ), .A3(_05102_ ), .ZN(_05103_ ) );
AOI211_X1 _12519_ ( .A(_04460_ ), .B(_05078_ ), .C1(_05084_ ), .C2(_05103_ ), .ZN(_00319_ ) );
XNOR2_X1 _12520_ ( .A(_05079_ ), .B(_03241_ ), .ZN(_05104_ ) );
NAND2_X1 _12521_ ( .A1(_05104_ ), .A2(_04550_ ), .ZN(_05105_ ) );
NAND3_X1 _12522_ ( .A1(_04889_ ), .A2(_04890_ ), .A3(_04508_ ), .ZN(_05106_ ) );
OR2_X1 _12523_ ( .A1(_04896_ ), .A2(_04865_ ), .ZN(_05107_ ) );
AND3_X1 _12524_ ( .A1(_05106_ ), .A2(_04757_ ), .A3(_05107_ ), .ZN(_05108_ ) );
AND2_X1 _12525_ ( .A1(_03475_ ), .A2(_04507_ ), .ZN(_05109_ ) );
AND3_X1 _12526_ ( .A1(\u_exu.alu_p1 [31] ), .A2(\u_exu.alu_ctrl [1] ), .A3(\u_exu.alu_p2 [3] ), .ZN(_05110_ ) );
OAI21_X1 _12527_ ( .A(\u_exu.alu_p2 [4] ), .B1(_05109_ ), .B2(_05110_ ), .ZN(_05111_ ) );
AND3_X1 _12528_ ( .A1(_03447_ ), .A2(_03455_ ), .A3(\u_exu.alu_p2 [3] ), .ZN(_05112_ ) );
AOI21_X1 _12529_ ( .A(\u_exu.alu_p2 [3] ), .B1(_03425_ ), .B2(_03432_ ), .ZN(_05113_ ) );
OAI21_X1 _12530_ ( .A(_04917_ ), .B1(_05112_ ), .B2(_05113_ ), .ZN(_05114_ ) );
AOI21_X1 _12531_ ( .A(_03437_ ), .B1(_05111_ ), .B2(_05114_ ), .ZN(_05115_ ) );
AOI211_X1 _12532_ ( .A(_05108_ ), .B(_05115_ ), .C1(_03117_ ), .C2(_04767_ ), .ZN(_05116_ ) );
AOI21_X1 _12533_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [8] ), .B2(\u_exu.alu_p2 [8] ), .ZN(_05117_ ) );
OAI211_X1 _12534_ ( .A(_04982_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [8] ), .C2(\u_exu.alu_p2 [8] ), .ZN(_05118_ ) );
OAI211_X1 _12535_ ( .A(_05105_ ), .B(_05116_ ), .C1(_05117_ ), .C2(_05118_ ), .ZN(_05119_ ) );
MUX2_X1 _12536_ ( .A(\u_exu.alu_p1 [8] ), .B(_05119_ ), .S(_04900_ ), .Z(_05120_ ) );
AND2_X1 _12537_ ( .A1(_05120_ ), .A2(_04593_ ), .ZN(_00320_ ) );
AOI21_X1 _12538_ ( .A(_03261_ ), .B1(_03277_ ), .B2(_03281_ ), .ZN(_05121_ ) );
INV_X1 _12539_ ( .A(_03288_ ), .ZN(_05122_ ) );
OAI21_X1 _12540_ ( .A(_03247_ ), .B1(_05121_ ), .B2(_05122_ ), .ZN(_05123_ ) );
NAND2_X1 _12541_ ( .A1(_03245_ ), .A2(\u_exu.alu_p1 [6] ), .ZN(_05124_ ) );
AND3_X1 _12542_ ( .A1(_05123_ ), .A2(_03250_ ), .A3(_05124_ ), .ZN(_05125_ ) );
AOI21_X1 _12543_ ( .A(_03250_ ), .B1(_05123_ ), .B2(_05124_ ), .ZN(_05126_ ) );
OAI21_X1 _12544_ ( .A(_04550_ ), .B1(_05125_ ), .B2(_05126_ ), .ZN(_05127_ ) );
NOR4_X1 _12545_ ( .A1(_03131_ ), .A2(_04723_ ), .A3(_04486_ ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_05128_ ) );
OAI21_X1 _12546_ ( .A(_05128_ ), .B1(fanout_net_11 ), .B2(_03130_ ), .ZN(_05129_ ) );
OAI21_X1 _12547_ ( .A(_04536_ ), .B1(_04538_ ), .B2(_04544_ ), .ZN(_05130_ ) );
AND3_X1 _12548_ ( .A1(_05130_ ), .A2(_04508_ ), .A3(_04756_ ), .ZN(_05131_ ) );
AND2_X1 _12549_ ( .A1(_04919_ ), .A2(_04865_ ), .ZN(_05132_ ) );
NOR3_X1 _12550_ ( .A1(_04929_ ), .A2(\u_exu.alu_ctrl [1] ), .A3(_04629_ ), .ZN(_05133_ ) );
NOR4_X1 _12551_ ( .A1(_05132_ ), .A2(_04917_ ), .A3(_05110_ ), .A4(_05133_ ), .ZN(_05134_ ) );
NAND3_X1 _12552_ ( .A1(_04924_ ), .A2(_04926_ ), .A3(\u_exu.alu_p2 [3] ), .ZN(_05135_ ) );
NAND3_X1 _12553_ ( .A1(_05045_ ), .A2(fanout_net_17 ), .A3(_05046_ ), .ZN(_05136_ ) );
OR3_X1 _12554_ ( .A1(_04529_ ), .A2(\u_exu.alu_p2 [1] ), .A3(_04518_ ), .ZN(_05137_ ) );
OR3_X1 _12555_ ( .A1(_04517_ ), .A2(_04527_ ), .A3(_04522_ ), .ZN(_05138_ ) );
AND2_X1 _12556_ ( .A1(_05137_ ), .A2(_05138_ ), .ZN(_05139_ ) );
OAI211_X1 _12557_ ( .A(_05136_ ), .B(_04507_ ), .C1(_05139_ ), .C2(fanout_net_17 ), .ZN(_05140_ ) );
AND3_X1 _12558_ ( .A1(_05135_ ), .A2(_05140_ ), .A3(_04618_ ), .ZN(_05141_ ) );
NOR3_X1 _12559_ ( .A1(_05134_ ), .A2(_03437_ ), .A3(_05141_ ), .ZN(_05142_ ) );
AOI211_X1 _12560_ ( .A(_05131_ ), .B(_05142_ ), .C1(_03132_ ), .C2(_04767_ ), .ZN(_05143_ ) );
NAND4_X1 _12561_ ( .A1(_05127_ ), .A2(_04879_ ), .A3(_05129_ ), .A4(_05143_ ), .ZN(_05144_ ) );
OAI21_X1 _12562_ ( .A(_05144_ ), .B1(\u_exu.alu_p1 [7] ), .B2(_04900_ ), .ZN(_05145_ ) );
NOR2_X1 _12563_ ( .A1(_05145_ ), .A2(_04472_ ), .ZN(_00321_ ) );
OAI21_X1 _12564_ ( .A(_04640_ ), .B1(_04643_ ), .B2(_04537_ ), .ZN(_05146_ ) );
AND3_X1 _12565_ ( .A1(_05146_ ), .A2(_04869_ ), .A3(_04588_ ), .ZN(_05147_ ) );
NOR2_X1 _12566_ ( .A1(_04944_ ), .A2(\u_exu.alu_p2 [3] ), .ZN(_05148_ ) );
NOR4_X1 _12567_ ( .A1(_03460_ ), .A2(_03099_ ), .A3(fanout_net_17 ), .A4(\u_exu.alu_p2 [1] ), .ZN(_05149_ ) );
OAI21_X1 _12568_ ( .A(_04930_ ), .B1(_05148_ ), .B2(_05149_ ), .ZN(_05150_ ) );
AOI21_X1 _12569_ ( .A(_04493_ ), .B1(_04600_ ), .B2(_04601_ ), .ZN(_05151_ ) );
OAI21_X1 _12570_ ( .A(_04605_ ), .B1(_05148_ ), .B2(_05151_ ), .ZN(_05152_ ) );
AOI21_X1 _12571_ ( .A(_04494_ ), .B1(_05062_ ), .B2(_05063_ ), .ZN(_05153_ ) );
OAI21_X1 _12572_ ( .A(_04527_ ), .B1(_03414_ ), .B2(_03415_ ), .ZN(_05154_ ) );
OAI21_X1 _12573_ ( .A(\u_exu.alu_p2 [1] ), .B1(_03422_ ), .B2(_03423_ ), .ZN(_05155_ ) );
AND2_X1 _12574_ ( .A1(_05154_ ), .A2(_05155_ ), .ZN(_05156_ ) );
AOI211_X1 _12575_ ( .A(\u_exu.alu_p2 [3] ), .B(_05153_ ), .C1(_04537_ ), .C2(_05156_ ), .ZN(_05157_ ) );
AOI21_X1 _12576_ ( .A(_05157_ ), .B1(\u_exu.alu_p2 [3] ), .B2(_04950_ ), .ZN(_05158_ ) );
OAI211_X1 _12577_ ( .A(_05150_ ), .B(_05152_ ), .C1(\u_exu.alu_p2 [4] ), .C2(_05158_ ), .ZN(_05159_ ) );
AOI221_X4 _12578_ ( .A(_05147_ ), .B1(_03107_ ), .B2(_03482_ ), .C1(_05159_ ), .C2(_04737_ ), .ZN(_05160_ ) );
OR3_X1 _12579_ ( .A1(_05121_ ), .A2(_03247_ ), .A3(_05122_ ), .ZN(_05161_ ) );
NAND3_X1 _12580_ ( .A1(_05161_ ), .A2(_04549_ ), .A3(_05123_ ), .ZN(_05162_ ) );
AOI21_X1 _12581_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [6] ), .B2(\u_exu.alu_p2 [6] ), .ZN(_05163_ ) );
OAI211_X1 _12582_ ( .A(_04982_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [6] ), .C2(\u_exu.alu_p2 [6] ), .ZN(_05164_ ) );
OAI211_X1 _12583_ ( .A(_05160_ ), .B(_05162_ ), .C1(_05163_ ), .C2(_05164_ ), .ZN(_05165_ ) );
MUX2_X1 _12584_ ( .A(\u_exu.alu_p1 [6] ), .B(_05165_ ), .S(_04879_ ), .Z(_05166_ ) );
AND2_X1 _12585_ ( .A1(_05166_ ), .A2(_04593_ ), .ZN(_00322_ ) );
AND2_X1 _12586_ ( .A1(_03277_ ), .A2(_03281_ ), .ZN(_05167_ ) );
INV_X1 _12587_ ( .A(_03256_ ), .ZN(_05168_ ) );
OR2_X1 _12588_ ( .A1(_05167_ ), .A2(_05168_ ), .ZN(_05169_ ) );
INV_X1 _12589_ ( .A(_03287_ ), .ZN(_05170_ ) );
AND3_X1 _12590_ ( .A1(_05169_ ), .A2(_03259_ ), .A3(_05170_ ), .ZN(_05171_ ) );
AOI21_X1 _12591_ ( .A(_03259_ ), .B1(_05169_ ), .B2(_05170_ ), .ZN(_05172_ ) );
OAI21_X1 _12592_ ( .A(_04550_ ), .B1(_05171_ ), .B2(_05172_ ), .ZN(_05173_ ) );
AND3_X1 _12593_ ( .A1(_04714_ ), .A2(_04869_ ), .A3(_04756_ ), .ZN(_05174_ ) );
OAI21_X1 _12594_ ( .A(_04930_ ), .B1(_04671_ ), .B2(_04675_ ), .ZN(_05175_ ) );
AND3_X1 _12595_ ( .A1(_05090_ ), .A2(fanout_net_17 ), .A3(_05091_ ), .ZN(_05176_ ) );
OAI21_X1 _12596_ ( .A(_04528_ ), .B1(_04532_ ), .B2(_04530_ ), .ZN(_05177_ ) );
OAI21_X1 _12597_ ( .A(\u_exu.alu_p2 [1] ), .B1(_04529_ ), .B2(_04518_ ), .ZN(_05178_ ) );
AOI21_X1 _12598_ ( .A(fanout_net_17 ), .B1(_05177_ ), .B2(_05178_ ), .ZN(_05179_ ) );
NOR2_X1 _12599_ ( .A1(_05176_ ), .A2(_05179_ ), .ZN(_05180_ ) );
MUX2_X1 _12600_ ( .A(_05180_ ), .B(_04970_ ), .S(\u_exu.alu_p2 [3] ), .Z(_05181_ ) );
OAI221_X1 _12601_ ( .A(_05175_ ), .B1(_05181_ ), .B2(\u_exu.alu_p2 [4] ), .C1(_04940_ ), .C2(_04683_ ), .ZN(_05182_ ) );
AOI221_X4 _12602_ ( .A(_05174_ ), .B1(_03109_ ), .B2(_04646_ ), .C1(_05182_ ), .C2(_04737_ ), .ZN(_05183_ ) );
AOI21_X1 _12603_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p1 [5] ), .B2(\u_exu.alu_p2 [5] ), .ZN(_05184_ ) );
OAI211_X1 _12604_ ( .A(_04982_ ), .B(fanout_net_19 ), .C1(\u_exu.alu_p1 [5] ), .C2(\u_exu.alu_p2 [5] ), .ZN(_05185_ ) );
OAI211_X1 _12605_ ( .A(_05173_ ), .B(_05183_ ), .C1(_05184_ ), .C2(_05185_ ), .ZN(_05186_ ) );
MUX2_X1 _12606_ ( .A(\u_exu.alu_p1 [5] ), .B(_05186_ ), .S(_04900_ ), .Z(_05187_ ) );
CLKBUF_X2 _12607_ ( .A(_04473_ ), .Z(_05188_ ) );
AND2_X1 _12608_ ( .A1(_05187_ ), .A2(_05188_ ), .ZN(_00323_ ) );
NAND3_X1 _12609_ ( .A1(_03277_ ), .A2(_03281_ ), .A3(_05168_ ), .ZN(_05189_ ) );
NAND3_X1 _12610_ ( .A1(_05169_ ), .A2(_04549_ ), .A3(_05189_ ), .ZN(_05190_ ) );
NAND3_X1 _12611_ ( .A1(_03421_ ), .A2(_03424_ ), .A3(fanout_net_17 ), .ZN(_05191_ ) );
OAI211_X1 _12612_ ( .A(_05191_ ), .B(_04493_ ), .C1(fanout_net_17 ), .C2(_03417_ ), .ZN(_05192_ ) );
OAI21_X1 _12613_ ( .A(_05192_ ), .B1(_04998_ ), .B2(_04629_ ), .ZN(_05193_ ) );
OAI22_X1 _12614_ ( .A1(_04735_ ), .A2(_04940_ ), .B1(\u_exu.alu_p2 [4] ), .B2(_05193_ ), .ZN(_05194_ ) );
NOR2_X1 _12615_ ( .A1(_04731_ ), .A2(_04931_ ), .ZN(_05195_ ) );
OAI21_X1 _12616_ ( .A(_04686_ ), .B1(_05194_ ), .B2(_05195_ ), .ZN(_05196_ ) );
NAND3_X1 _12617_ ( .A1(_04762_ ), .A2(_04508_ ), .A3(_04756_ ), .ZN(_05197_ ) );
AND2_X1 _12618_ ( .A1(_05196_ ), .A2(_05197_ ), .ZN(_05198_ ) );
AOI21_X1 _12619_ ( .A(_03481_ ), .B1(_04917_ ), .B2(_03255_ ), .ZN(_05199_ ) );
AND2_X1 _12620_ ( .A1(\u_exu.alu_p2 [4] ), .A2(\u_exu.alu_p1 [4] ), .ZN(_05200_ ) );
OAI21_X1 _12621_ ( .A(_05199_ ), .B1(fanout_net_11 ), .B2(_05200_ ), .ZN(_05201_ ) );
NAND2_X1 _12622_ ( .A1(_03127_ ), .A2(_04646_ ), .ZN(_05202_ ) );
NAND4_X1 _12623_ ( .A1(_05190_ ), .A2(_05198_ ), .A3(_05201_ ), .A4(_05202_ ), .ZN(_05203_ ) );
MUX2_X1 _12624_ ( .A(\u_exu.alu_p1 [4] ), .B(_05203_ ), .S(_04653_ ), .Z(_05204_ ) );
AND2_X1 _12625_ ( .A1(_05204_ ), .A2(_05188_ ), .ZN(_00324_ ) );
AND4_X1 _12626_ ( .A1(\u_exu.alu_p1 [3] ), .A2(_04486_ ), .A3(_04487_ ), .A4(fanout_net_19 ), .ZN(_05205_ ) );
NOR2_X1 _12627_ ( .A1(_03274_ ), .A2(_03276_ ), .ZN(_05206_ ) );
NOR2_X1 _12628_ ( .A1(_03266_ ), .A2(\u_exu.alu_p1 [2] ), .ZN(_05207_ ) );
NOR3_X1 _12629_ ( .A1(_05206_ ), .A2(_03278_ ), .A3(_05207_ ), .ZN(_05208_ ) );
OR3_X1 _12630_ ( .A1(_05208_ ), .A2(_03264_ ), .A3(_03278_ ), .ZN(_05209_ ) );
OAI21_X1 _12631_ ( .A(_03264_ ), .B1(_05208_ ), .B2(_03278_ ), .ZN(_05210_ ) );
AND3_X1 _12632_ ( .A1(_05209_ ), .A2(_04549_ ), .A3(_05210_ ), .ZN(_05211_ ) );
OAI211_X1 _12633_ ( .A(_04649_ ), .B(fanout_net_19 ), .C1(fanout_net_11 ), .C2(\u_exu.alu_p1 [3] ), .ZN(_05212_ ) );
NAND2_X1 _12634_ ( .A1(fanout_net_11 ), .A2(\u_exu.alu_p1 [3] ), .ZN(_05213_ ) );
AOI21_X1 _12635_ ( .A(_05212_ ), .B1(_04754_ ), .B2(_05213_ ), .ZN(_05214_ ) );
AND2_X1 _12636_ ( .A1(_03108_ ), .A2(_04646_ ), .ZN(_05215_ ) );
OAI21_X1 _12637_ ( .A(_04605_ ), .B1(_04790_ ), .B2(_04786_ ), .ZN(_05216_ ) );
OAI21_X1 _12638_ ( .A(_04930_ ), .B1(_04779_ ), .B2(_04786_ ), .ZN(_05217_ ) );
OAI21_X1 _12639_ ( .A(\u_exu.alu_p2 [1] ), .B1(_04532_ ), .B2(_04530_ ), .ZN(_05218_ ) );
NOR2_X1 _12640_ ( .A1(_04539_ ), .A2(_04533_ ), .ZN(_05219_ ) );
OAI211_X1 _12641_ ( .A(_05218_ ), .B(_04494_ ), .C1(_05219_ ), .C2(\u_exu.alu_p2 [1] ), .ZN(_05220_ ) );
OAI21_X1 _12642_ ( .A(_05220_ ), .B1(_04495_ ), .B2(_05139_ ), .ZN(_05221_ ) );
MUX2_X1 _12643_ ( .A(_05048_ ), .B(_05221_ ), .S(_04629_ ), .Z(_05222_ ) );
OAI211_X1 _12644_ ( .A(_05216_ ), .B(_05217_ ), .C1(_05222_ ), .C2(\u_exu.alu_p2 [4] ), .ZN(_05223_ ) );
NAND2_X1 _12645_ ( .A1(_05223_ ), .A2(_04686_ ), .ZN(_05224_ ) );
NAND3_X1 _12646_ ( .A1(_04793_ ), .A2(_04508_ ), .A3(_04756_ ), .ZN(_05225_ ) );
NAND2_X1 _12647_ ( .A1(_05224_ ), .A2(_05225_ ), .ZN(_05226_ ) );
OR4_X1 _12648_ ( .A1(_05211_ ), .A2(_05214_ ), .A3(_05215_ ), .A4(_05226_ ), .ZN(_05227_ ) );
AOI21_X1 _12649_ ( .A(_05205_ ), .B1(_05227_ ), .B2(_04900_ ), .ZN(_05228_ ) );
NOR2_X1 _12650_ ( .A1(_05228_ ), .A2(_04472_ ), .ZN(_00325_ ) );
AND4_X1 _12651_ ( .A1(_04618_ ), .A2(_04808_ ), .A3(_04865_ ), .A4(_03104_ ), .ZN(_05229_ ) );
NOR2_X1 _12652_ ( .A1(_03411_ ), .A2(_03412_ ), .ZN(_05230_ ) );
MUX2_X1 _12653_ ( .A(_05230_ ), .B(_03407_ ), .S(_04527_ ), .Z(_05231_ ) );
MUX2_X1 _12654_ ( .A(_05156_ ), .B(_05231_ ), .S(_04494_ ), .Z(_05232_ ) );
AOI21_X1 _12655_ ( .A(\u_exu.alu_p2 [4] ), .B1(_05232_ ), .B2(_04507_ ), .ZN(_05233_ ) );
OAI21_X1 _12656_ ( .A(_05233_ ), .B1(_04869_ ), .B2(_05066_ ), .ZN(_05234_ ) );
OAI221_X1 _12657_ ( .A(_05234_ ), .B1(_04827_ ), .B2(_04931_ ), .C1(_04830_ ), .C2(_04940_ ), .ZN(_05235_ ) );
AOI221_X4 _12658_ ( .A(_05229_ ), .B1(_03129_ ), .B2(_04646_ ), .C1(_05235_ ), .C2(_04737_ ), .ZN(_05236_ ) );
XNOR2_X1 _12659_ ( .A(_05206_ ), .B(_03268_ ), .ZN(_05237_ ) );
NAND2_X1 _12660_ ( .A1(_05237_ ), .A2(_04550_ ), .ZN(_05238_ ) );
AOI21_X1 _12661_ ( .A(fanout_net_11 ), .B1(fanout_net_17 ), .B2(\u_exu.alu_p1 [2] ), .ZN(_05239_ ) );
OAI211_X1 _12662_ ( .A(_04982_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p2 [2] ), .C2(\u_exu.alu_p1 [2] ), .ZN(_05240_ ) );
OAI211_X1 _12663_ ( .A(_05236_ ), .B(_05238_ ), .C1(_05239_ ), .C2(_05240_ ), .ZN(_05241_ ) );
MUX2_X1 _12664_ ( .A(\u_exu.alu_p1 [2] ), .B(_05241_ ), .S(_04879_ ), .Z(_05242_ ) );
AND2_X1 _12665_ ( .A1(_05242_ ), .A2(_05188_ ), .ZN(_00326_ ) );
NOR4_X1 _12666_ ( .A1(_05007_ ), .A2(_04723_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03490_ ), .ZN(_05243_ ) );
NAND3_X1 _12667_ ( .A1(_03369_ ), .A2(_03381_ ), .A3(_03184_ ), .ZN(_05244_ ) );
NAND2_X1 _12668_ ( .A1(_05243_ ), .A2(_05244_ ), .ZN(_05245_ ) );
NOR4_X1 _12669_ ( .A1(_03144_ ), .A2(_04723_ ), .A3(_03400_ ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_05246_ ) );
OAI21_X1 _12670_ ( .A(_05246_ ), .B1(fanout_net_11 ), .B2(_03143_ ), .ZN(_05247_ ) );
NAND3_X1 _12671_ ( .A1(_03145_ ), .A2(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .A3(_03092_ ), .ZN(_05248_ ) );
AND2_X1 _12672_ ( .A1(_04993_ ), .A2(_04865_ ), .ZN(_05249_ ) );
OAI21_X1 _12673_ ( .A(_04977_ ), .B1(_05249_ ), .B2(\u_exu.alu_ctrl [1] ), .ZN(_05250_ ) );
OR2_X1 _12674_ ( .A1(_05000_ ), .A2(\u_exu.alu_p2 [4] ), .ZN(_05251_ ) );
AND2_X1 _12675_ ( .A1(\u_exu.alu_p1 [31] ), .A2(\u_exu.alu_p2 [4] ), .ZN(_05252_ ) );
INV_X1 _12676_ ( .A(_05252_ ), .ZN(_05253_ ) );
AOI21_X1 _12677_ ( .A(_05250_ ), .B1(_05251_ ), .B2(_05253_ ), .ZN(_05254_ ) );
OAI211_X1 _12678_ ( .A(_03466_ ), .B(_04491_ ), .C1(\u_exu.alu_p2 [0] ), .C2(_03182_ ), .ZN(_05255_ ) );
NAND3_X1 _12679_ ( .A1(_03464_ ), .A2(\u_exu.alu_p2 [1] ), .A3(_03472_ ), .ZN(_05256_ ) );
NAND3_X1 _12680_ ( .A1(_05255_ ), .A2(_05256_ ), .A3(_04495_ ), .ZN(_05257_ ) );
NOR2_X1 _12681_ ( .A1(_04620_ ), .A2(_03449_ ), .ZN(_05258_ ) );
MUX2_X1 _12682_ ( .A(_05258_ ), .B(_04615_ ), .S(_04528_ ), .Z(_05259_ ) );
OAI211_X1 _12683_ ( .A(_04507_ ), .B(_05257_ ), .C1(_05259_ ), .C2(_04516_ ), .ZN(_05260_ ) );
NAND3_X1 _12684_ ( .A1(_04750_ ), .A2(_04753_ ), .A3(\u_exu.alu_p2 [3] ), .ZN(_05261_ ) );
AND3_X1 _12685_ ( .A1(_05260_ ), .A2(_04618_ ), .A3(_05261_ ), .ZN(_05262_ ) );
AND2_X1 _12686_ ( .A1(_05262_ ), .A2(_03104_ ), .ZN(_05263_ ) );
INV_X1 _12687_ ( .A(_04506_ ), .ZN(_05264_ ) );
NOR2_X1 _12688_ ( .A1(_04991_ ), .A2(_05264_ ), .ZN(_05265_ ) );
NOR3_X1 _12689_ ( .A1(_05254_ ), .A2(_05263_ ), .A3(_05265_ ), .ZN(_05266_ ) );
NAND4_X1 _12690_ ( .A1(_05245_ ), .A2(_05247_ ), .A3(_05248_ ), .A4(_05266_ ), .ZN(_05267_ ) );
MUX2_X1 _12691_ ( .A(\u_exu.alu_p1 [28] ), .B(_05267_ ), .S(_04879_ ), .Z(_05268_ ) );
AND2_X1 _12692_ ( .A1(_05268_ ), .A2(_05188_ ), .ZN(_00327_ ) );
AND4_X1 _12693_ ( .A1(_04618_ ), .A2(_04872_ ), .A3(_04869_ ), .A4(_03104_ ), .ZN(_05269_ ) );
OAI21_X1 _12694_ ( .A(_04605_ ), .B1(_04860_ ), .B2(_04855_ ), .ZN(_05270_ ) );
OAI21_X1 _12695_ ( .A(_04930_ ), .B1(_04850_ ), .B2(_04855_ ), .ZN(_05271_ ) );
AND2_X1 _12696_ ( .A1(_05177_ ), .A2(_05178_ ), .ZN(_05272_ ) );
MUX2_X1 _12697_ ( .A(_04542_ ), .B(_03267_ ), .S(\u_exu.alu_p2 [0] ), .Z(_05273_ ) );
MUX2_X1 _12698_ ( .A(_05273_ ), .B(_05219_ ), .S(\u_exu.alu_p2 [1] ), .Z(_05274_ ) );
MUX2_X1 _12699_ ( .A(_05272_ ), .B(_05274_ ), .S(_03102_ ), .Z(_05275_ ) );
AND2_X1 _12700_ ( .A1(_05275_ ), .A2(_04869_ ), .ZN(_05276_ ) );
OAI21_X1 _12701_ ( .A(_04618_ ), .B1(_05093_ ), .B2(_04869_ ), .ZN(_05277_ ) );
OAI211_X1 _12702_ ( .A(_05270_ ), .B(_05271_ ), .C1(_05276_ ), .C2(_05277_ ), .ZN(_05278_ ) );
AOI221_X4 _12703_ ( .A(_05269_ ), .B1(_03128_ ), .B2(_04646_ ), .C1(_05278_ ), .C2(_04737_ ), .ZN(_05279_ ) );
NOR4_X1 _12704_ ( .A1(_03274_ ), .A2(_04724_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_04487_ ), .ZN(_05280_ ) );
AOI21_X1 _12705_ ( .A(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .B1(_03084_ ), .B2(\u_exu.alu_p2 [0] ), .ZN(_05281_ ) );
NOR3_X1 _12706_ ( .A1(_03089_ ), .A2(\u_exu.alu_ctrl [3] ), .A3(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ), .ZN(_05282_ ) );
OR3_X1 _12707_ ( .A1(_03271_ ), .A2(_05281_ ), .A3(_05282_ ), .ZN(_05283_ ) );
NAND2_X1 _12708_ ( .A1(_05280_ ), .A2(_05283_ ), .ZN(_05284_ ) );
OAI211_X1 _12709_ ( .A(_04649_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p2 [1] ), .C2(\u_exu.alu_p1 [1] ), .ZN(_05285_ ) );
AOI21_X1 _12710_ ( .A(fanout_net_11 ), .B1(\u_exu.alu_p2 [1] ), .B2(\u_exu.alu_p1 [1] ), .ZN(_05286_ ) );
OR2_X1 _12711_ ( .A1(_05285_ ), .A2(_05286_ ), .ZN(_05287_ ) );
AND4_X1 _12712_ ( .A1(_04879_ ), .A2(_05279_ ), .A3(_05284_ ), .A4(_05287_ ), .ZN(_05288_ ) );
AND4_X1 _12713_ ( .A1(_04542_ ), .A2(_04486_ ), .A3(_04487_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05289_ ) );
NOR3_X1 _12714_ ( .A1(_05288_ ), .A2(_04470_ ), .A3(_05289_ ), .ZN(_00328_ ) );
AND3_X1 _12715_ ( .A1(_03489_ ), .A2(_04476_ ), .A3(_03491_ ), .ZN(_00329_ ) );
INV_X1 _12716_ ( .A(_03360_ ), .ZN(_05290_ ) );
INV_X1 _12717_ ( .A(_03375_ ), .ZN(_05291_ ) );
INV_X1 _12718_ ( .A(_03365_ ), .ZN(_05292_ ) );
AOI21_X1 _12719_ ( .A(_05292_ ), .B1(_03327_ ), .B2(_03350_ ), .ZN(_05293_ ) );
OAI21_X1 _12720_ ( .A(_05291_ ), .B1(_05293_ ), .B2(_03373_ ), .ZN(_05294_ ) );
AOI21_X1 _12721_ ( .A(_05290_ ), .B1(_05294_ ), .B2(_03372_ ), .ZN(_05295_ ) );
OR3_X1 _12722_ ( .A1(_05295_ ), .A2(_03356_ ), .A3(_03379_ ), .ZN(_05296_ ) );
OAI21_X1 _12723_ ( .A(_03356_ ), .B1(_05295_ ), .B2(_03379_ ), .ZN(_05297_ ) );
NAND3_X1 _12724_ ( .A1(_05296_ ), .A2(_04550_ ), .A3(_05297_ ), .ZN(_05298_ ) );
AND2_X1 _12725_ ( .A1(_04580_ ), .A2(_04585_ ), .ZN(_05299_ ) );
MUX2_X1 _12726_ ( .A(_04566_ ), .B(_05299_ ), .S(\u_exu.alu_p2 [2] ), .Z(_05300_ ) );
MUX2_X1 _12727_ ( .A(_04804_ ), .B(_05300_ ), .S(_04493_ ), .Z(_05301_ ) );
NAND2_X1 _12728_ ( .A1(_05301_ ), .A2(_04756_ ), .ZN(_05302_ ) );
NAND3_X1 _12729_ ( .A1(_05037_ ), .A2(_05038_ ), .A3(_04505_ ), .ZN(_05303_ ) );
NAND2_X1 _12730_ ( .A1(_05302_ ), .A2(_05303_ ), .ZN(_05304_ ) );
OAI21_X1 _12731_ ( .A(_05253_ ), .B1(_05043_ ), .B2(\u_exu.alu_p2 [4] ), .ZN(_05305_ ) );
NAND2_X1 _12732_ ( .A1(_04778_ ), .A2(_04630_ ), .ZN(_05306_ ) );
AOI21_X1 _12733_ ( .A(_04978_ ), .B1(_05306_ ), .B2(_04497_ ), .ZN(_05307_ ) );
AOI221_X4 _12734_ ( .A(_05304_ ), .B1(_03122_ ), .B2(_04646_ ), .C1(_05305_ ), .C2(_05307_ ), .ZN(_05308_ ) );
AOI21_X1 _12735_ ( .A(\u_exu.alu_ctrl [0] ), .B1(\u_exu.alu_p1 [27] ), .B2(\u_exu.alu_p2 [27] ), .ZN(_05309_ ) );
OAI211_X1 _12736_ ( .A(_04982_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1 [27] ), .C2(\u_exu.alu_p2 [27] ), .ZN(_05310_ ) );
OAI211_X1 _12737_ ( .A(_05298_ ), .B(_05308_ ), .C1(_05309_ ), .C2(_05310_ ), .ZN(_05311_ ) );
MUX2_X1 _12738_ ( .A(\u_exu.alu_p1 [27] ), .B(_05311_ ), .S(_04879_ ), .Z(_05312_ ) );
AND2_X1 _12739_ ( .A1(_05312_ ), .A2(_05188_ ), .ZN(_00330_ ) );
NOR4_X1 _12740_ ( .A1(_05295_ ), .A2(_04724_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03490_ ), .ZN(_05313_ ) );
NAND3_X1 _12741_ ( .A1(_05294_ ), .A2(_05290_ ), .A3(_03372_ ), .ZN(_05314_ ) );
NAND2_X1 _12742_ ( .A1(_05313_ ), .A2(_05314_ ), .ZN(_05315_ ) );
OAI21_X1 _12743_ ( .A(_04917_ ), .B1(_05070_ ), .B2(_04603_ ), .ZN(_05316_ ) );
AOI21_X1 _12744_ ( .A(_04497_ ), .B1(_05316_ ), .B2(_05253_ ), .ZN(_05317_ ) );
AND4_X1 _12745_ ( .A1(_04497_ ), .A2(_04825_ ), .A3(_04618_ ), .A4(_04869_ ), .ZN(_05318_ ) );
OAI21_X1 _12746_ ( .A(_04737_ ), .B1(_05317_ ), .B2(_05318_ ), .ZN(_05319_ ) );
NAND3_X1 _12747_ ( .A1(_05059_ ), .A2(_05060_ ), .A3(_04506_ ), .ZN(_05320_ ) );
NAND3_X1 _12748_ ( .A1(_04619_ ), .A2(_04621_ ), .A3(\u_exu.alu_p2 [2] ), .ZN(_05321_ ) );
OAI211_X1 _12749_ ( .A(_05321_ ), .B(_04508_ ), .C1(_04616_ ), .C2(\u_exu.alu_p2 [2] ), .ZN(_05322_ ) );
NAND3_X1 _12750_ ( .A1(_04839_ ), .A2(_04840_ ), .A3(\u_exu.alu_p2 [3] ), .ZN(_05323_ ) );
NAND3_X1 _12751_ ( .A1(_05322_ ), .A2(_04757_ ), .A3(_05323_ ), .ZN(_05324_ ) );
NAND2_X1 _12752_ ( .A1(_03141_ ), .A2(_04767_ ), .ZN(_05325_ ) );
AND4_X1 _12753_ ( .A1(_05319_ ), .A2(_05320_ ), .A3(_05324_ ), .A4(_05325_ ), .ZN(_05326_ ) );
AOI21_X1 _12754_ ( .A(\u_exu.alu_ctrl [0] ), .B1(\u_exu.alu_p1 [26] ), .B2(\u_exu.alu_p2 [26] ), .ZN(_05327_ ) );
OAI211_X1 _12755_ ( .A(_04982_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1 [26] ), .C2(\u_exu.alu_p2 [26] ), .ZN(_05328_ ) );
OAI211_X1 _12756_ ( .A(_05315_ ), .B(_05326_ ), .C1(_05327_ ), .C2(_05328_ ), .ZN(_05329_ ) );
MUX2_X1 _12757_ ( .A(\u_exu.alu_p1 [26] ), .B(_05329_ ), .S(_04900_ ), .Z(_05330_ ) );
AND2_X1 _12758_ ( .A1(_05330_ ), .A2(_05188_ ), .ZN(_00331_ ) );
AND4_X1 _12759_ ( .A1(_03370_ ), .A2(_04486_ ), .A3(_04487_ ), .A4(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .ZN(_05331_ ) );
OR3_X1 _12760_ ( .A1(_05293_ ), .A2(_03373_ ), .A3(_03368_ ), .ZN(_05332_ ) );
OAI21_X1 _12761_ ( .A(_03368_ ), .B1(_05293_ ), .B2(_03373_ ), .ZN(_05333_ ) );
NAND3_X1 _12762_ ( .A1(_05332_ ), .A2(_04550_ ), .A3(_05333_ ), .ZN(_05334_ ) );
AOI21_X1 _12763_ ( .A(_05264_ ), .B1(_05085_ ), .B2(_05086_ ), .ZN(_05335_ ) );
AND3_X1 _12764_ ( .A1(_05020_ ), .A2(_05021_ ), .A3(_04537_ ), .ZN(_05336_ ) );
AOI211_X1 _12765_ ( .A(\u_exu.alu_p2 [3] ), .B(_05336_ ), .C1(\u_exu.alu_p2 [2] ), .C2(_04690_ ), .ZN(_05337_ ) );
AND3_X1 _12766_ ( .A1(_04863_ ), .A2(_04864_ ), .A3(\u_exu.alu_p2 [3] ), .ZN(_05338_ ) );
NOR3_X1 _12767_ ( .A1(_05337_ ), .A2(_04589_ ), .A3(_05338_ ), .ZN(_05339_ ) );
OAI21_X1 _12768_ ( .A(_05253_ ), .B1(_05098_ ), .B2(\u_exu.alu_p2 [4] ), .ZN(_05340_ ) );
AOI21_X1 _12769_ ( .A(_04978_ ), .B1(_05096_ ), .B2(_04497_ ), .ZN(_05341_ ) );
AOI211_X1 _12770_ ( .A(_05335_ ), .B(_05339_ ), .C1(_05340_ ), .C2(_05341_ ), .ZN(_05342_ ) );
NOR4_X1 _12771_ ( .A1(_03147_ ), .A2(_04723_ ), .A3(_03400_ ), .A4(\u_exu.alu_ctrl [4] ), .ZN(_05343_ ) );
OAI21_X1 _12772_ ( .A(_05343_ ), .B1(\u_exu.alu_ctrl [0] ), .B2(_03146_ ), .ZN(_05344_ ) );
NAND3_X1 _12773_ ( .A1(_03148_ ), .A2(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .A3(_03092_ ), .ZN(_05345_ ) );
AND4_X1 _12774_ ( .A1(_04653_ ), .A2(_05342_ ), .A3(_05344_ ), .A4(_05345_ ), .ZN(_05346_ ) );
AOI211_X1 _12775_ ( .A(_04460_ ), .B(_05331_ ), .C1(_05334_ ), .C2(_05346_ ), .ZN(_00332_ ) );
NOR4_X1 _12776_ ( .A1(_05293_ ), .A2(_04723_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03490_ ), .ZN(_05347_ ) );
OAI21_X1 _12777_ ( .A(_05347_ ), .B1(_03352_ ), .B2(_03365_ ), .ZN(_05348_ ) );
OAI21_X1 _12778_ ( .A(_04917_ ), .B1(_05109_ ), .B2(_04603_ ), .ZN(_05349_ ) );
AOI21_X1 _12779_ ( .A(_04497_ ), .B1(_05349_ ), .B2(_05253_ ), .ZN(_05350_ ) );
AND4_X1 _12780_ ( .A1(_04497_ ), .A2(_03475_ ), .A3(_04618_ ), .A4(_04869_ ), .ZN(_05351_ ) );
OAI21_X1 _12781_ ( .A(_04737_ ), .B1(_05350_ ), .B2(_05351_ ), .ZN(_05352_ ) );
NAND3_X1 _12782_ ( .A1(_05106_ ), .A2(_04506_ ), .A3(_05107_ ), .ZN(_05353_ ) );
AOI21_X1 _12783_ ( .A(_04516_ ), .B1(_04751_ ), .B2(_04752_ ), .ZN(_05354_ ) );
AOI211_X1 _12784_ ( .A(\u_exu.alu_p2 [3] ), .B(_05354_ ), .C1(_04538_ ), .C2(_05259_ ), .ZN(_05355_ ) );
AOI21_X1 _12785_ ( .A(_04508_ ), .B1(_04892_ ), .B2(_04893_ ), .ZN(_05356_ ) );
OAI21_X1 _12786_ ( .A(_04757_ ), .B1(_05355_ ), .B2(_05356_ ), .ZN(_05357_ ) );
NAND2_X1 _12787_ ( .A1(_04767_ ), .A2(_03124_ ), .ZN(_05358_ ) );
AND4_X1 _12788_ ( .A1(_05352_ ), .A2(_05353_ ), .A3(_05357_ ), .A4(_05358_ ), .ZN(_05359_ ) );
AOI21_X1 _12789_ ( .A(\u_exu.alu_ctrl [0] ), .B1(\u_exu.alu_p1 [24] ), .B2(\u_exu.alu_p2 [24] ), .ZN(_05360_ ) );
OAI211_X1 _12790_ ( .A(_04982_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1 [24] ), .C2(\u_exu.alu_p2 [24] ), .ZN(_05361_ ) );
OAI211_X1 _12791_ ( .A(_05348_ ), .B(_05359_ ), .C1(_05360_ ), .C2(_05361_ ), .ZN(_05362_ ) );
MUX2_X1 _12792_ ( .A(\u_exu.alu_p1 [24] ), .B(_05362_ ), .S(_04900_ ), .Z(_05363_ ) );
AND2_X1 _12793_ ( .A1(_05363_ ), .A2(_05188_ ), .ZN(_00333_ ) );
INV_X1 _12794_ ( .A(_03300_ ), .ZN(_05364_ ) );
NAND2_X1 _12795_ ( .A1(_04726_ ), .A2(_03309_ ), .ZN(_05365_ ) );
AOI21_X1 _12796_ ( .A(_05364_ ), .B1(_05365_ ), .B2(_03345_ ), .ZN(_05366_ ) );
OR3_X2 _12797_ ( .A1(_05366_ ), .A2(_03296_ ), .A3(_03348_ ), .ZN(_05367_ ) );
OAI21_X1 _12798_ ( .A(_03296_ ), .B1(_05366_ ), .B2(_03348_ ), .ZN(_05368_ ) );
AND3_X2 _12799_ ( .A1(_05367_ ), .A2(_04549_ ), .A3(_05368_ ), .ZN(_05369_ ) );
OAI21_X1 _12800_ ( .A(_04917_ ), .B1(_05132_ ), .B2(_05133_ ), .ZN(_05370_ ) );
OAI211_X1 _12801_ ( .A(\u_exu.alu_p1 [31] ), .B(\u_exu.alu_ctrl [1] ), .C1(\u_exu.alu_p2 [4] ), .C2(\u_exu.alu_p2 [3] ), .ZN(_05371_ ) );
AOI21_X1 _12802_ ( .A(_03437_ ), .B1(_05370_ ), .B2(_05371_ ), .ZN(_05372_ ) );
OAI21_X1 _12803_ ( .A(\u_exu.alu_p2 [3] ), .B1(_04515_ ), .B2(_04525_ ), .ZN(_05373_ ) );
NAND3_X1 _12804_ ( .A1(_04575_ ), .A2(_04586_ ), .A3(_04630_ ), .ZN(_05374_ ) );
AND3_X1 _12805_ ( .A1(_05373_ ), .A2(_04756_ ), .A3(_05374_ ), .ZN(_05375_ ) );
NAND3_X1 _12806_ ( .A1(_05130_ ), .A2(_04508_ ), .A3(_04506_ ), .ZN(_05376_ ) );
NAND2_X1 _12807_ ( .A1(_03111_ ), .A2(_03482_ ), .ZN(_05377_ ) );
AOI21_X1 _12808_ ( .A(\u_exu.alu_ctrl [0] ), .B1(\u_exu.alu_p1 [23] ), .B2(\u_exu.alu_p2 [23] ), .ZN(_05378_ ) );
OAI211_X1 _12809_ ( .A(_03401_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_p1 [23] ), .C2(\u_exu.alu_p2 [23] ), .ZN(_05379_ ) );
OAI211_X1 _12810_ ( .A(_05376_ ), .B(_05377_ ), .C1(_05378_ ), .C2(_05379_ ), .ZN(_05380_ ) );
OR4_X4 _12811_ ( .A1(_05369_ ), .A2(_05372_ ), .A3(_05375_ ), .A4(_05380_ ), .ZN(_05381_ ) );
MUX2_X2 _12812_ ( .A(\u_exu.alu_p1 [23] ), .B(_05381_ ), .S(_04879_ ), .Z(_05382_ ) );
AND2_X1 _12813_ ( .A1(_05382_ ), .A2(_05188_ ), .ZN(_00334_ ) );
NOR4_X1 _12814_ ( .A1(_05366_ ), .A2(_03435_ ), .A3(\u_exu.alu_ctrl [5] ), .A4(_03086_ ), .ZN(_05383_ ) );
NAND3_X1 _12815_ ( .A1(_05365_ ), .A2(_05364_ ), .A3(_03345_ ), .ZN(_05384_ ) );
NAND2_X1 _12816_ ( .A1(_05383_ ), .A2(_05384_ ), .ZN(_05385_ ) );
OAI21_X1 _12817_ ( .A(_04608_ ), .B1(_05148_ ), .B2(_05149_ ), .ZN(_05386_ ) );
OAI21_X1 _12818_ ( .A(_04599_ ), .B1(_05148_ ), .B2(_05151_ ), .ZN(_05387_ ) );
NAND2_X1 _12819_ ( .A1(_05386_ ), .A2(_05387_ ), .ZN(_05388_ ) );
OAI21_X1 _12820_ ( .A(_04686_ ), .B1(_05388_ ), .B2(_04606_ ), .ZN(_05389_ ) );
NOR3_X1 _12821_ ( .A1(_04633_ ), .A2(_04636_ ), .A3(_04865_ ), .ZN(_05390_ ) );
AOI21_X1 _12822_ ( .A(\u_exu.alu_p2 [3] ), .B1(_04622_ ), .B2(_04625_ ), .ZN(_05391_ ) );
OAI21_X1 _12823_ ( .A(_04756_ ), .B1(_05390_ ), .B2(_05391_ ), .ZN(_05392_ ) );
AND3_X1 _12824_ ( .A1(_05146_ ), .A2(_04865_ ), .A3(_04505_ ), .ZN(_05393_ ) );
OR4_X1 _12825_ ( .A1(_03435_ ), .A2(_03156_ ), .A3(_03400_ ), .A4(_03086_ ), .ZN(_05394_ ) );
OAI211_X1 _12826_ ( .A(_03401_ ), .B(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .C1(\u_exu.alu_ctrl [0] ), .C2(_03156_ ), .ZN(_05395_ ) );
AOI21_X1 _12827_ ( .A(_03157_ ), .B1(_05394_ ), .B2(_05395_ ), .ZN(_05396_ ) );
NOR2_X1 _12828_ ( .A1(_05393_ ), .A2(_05396_ ), .ZN(_05397_ ) );
NAND4_X1 _12829_ ( .A1(_05385_ ), .A2(_05389_ ), .A3(_05392_ ), .A4(_05397_ ), .ZN(_05398_ ) );
MUX2_X1 _12830_ ( .A(\u_exu.alu_p1 [22] ), .B(_05398_ ), .S(_04653_ ), .Z(_05399_ ) );
AND2_X1 _12831_ ( .A1(_05399_ ), .A2(_05188_ ), .ZN(_00335_ ) );
AOI21_X1 _12832_ ( .A(\u_ifu.jpc_ok_$_NOT__A_Y ), .B1(_00746_ ), .B2(_00758_ ), .ZN(_05400_ ) );
INV_X1 _12833_ ( .A(_00758_ ), .ZN(_05401_ ) );
AOI211_X1 _12834_ ( .A(idu_ready ), .B(_05401_ ), .C1(_00738_ ), .C2(_00745_ ), .ZN(_05402_ ) );
NOR2_X1 _12835_ ( .A1(_05400_ ), .A2(_05402_ ), .ZN(_05403_ ) );
INV_X1 _12836_ ( .A(_05403_ ), .ZN(_05404_ ) );
INV_X1 _12837_ ( .A(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ), .ZN(_05405_ ) );
INV_X1 _12838_ ( .A(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .ZN(_05406_ ) );
BUF_X4 _12839_ ( .A(_05406_ ), .Z(_05407_ ) );
NAND2_X1 _12840_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][23] ), .ZN(_05408_ ) );
NAND2_X1 _12841_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][23] ), .ZN(_05409_ ) );
AOI21_X1 _12842_ ( .A(\fc_addr [28] ), .B1(_05408_ ), .B2(_05409_ ), .ZN(_05410_ ) );
BUF_X4 _12843_ ( .A(_05407_ ), .Z(_05411_ ) );
NAND2_X1 _12844_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][25] ), .ZN(_05412_ ) );
NAND2_X1 _12845_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][25] ), .ZN(_05413_ ) );
AND3_X1 _12846_ ( .A1(_05412_ ), .A2(\fc_addr [30] ), .A3(_05413_ ), .ZN(_05414_ ) );
NOR2_X1 _12847_ ( .A1(_05411_ ), .A2(\u_icache.ctags[1][24] ), .ZN(_05415_ ) );
INV_X1 _12848_ ( .A(\fc_addr [29] ), .ZN(_05416_ ) );
NOR2_X1 _12849_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[0][24] ), .ZN(_05417_ ) );
OR3_X1 _12850_ ( .A1(_05415_ ), .A2(_05416_ ), .A3(_05417_ ), .ZN(_05418_ ) );
OAI21_X1 _12851_ ( .A(_05416_ ), .B1(_05415_ ), .B2(_05417_ ), .ZN(_05419_ ) );
AOI211_X1 _12852_ ( .A(_05410_ ), .B(_05414_ ), .C1(_05418_ ), .C2(_05419_ ), .ZN(_05420_ ) );
NAND2_X1 _12853_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][12] ), .ZN(_05421_ ) );
NAND2_X1 _12854_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][12] ), .ZN(_05422_ ) );
AND3_X1 _12855_ ( .A1(_05421_ ), .A2(\fc_addr [17] ), .A3(_05422_ ), .ZN(_05423_ ) );
MUX2_X1 _12856_ ( .A(\u_icache.ctags[0][8] ), .B(\u_icache.ctags[1][8] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05424_ ) );
INV_X1 _12857_ ( .A(\fc_addr [13] ), .ZN(_05425_ ) );
AND2_X1 _12858_ ( .A1(_05424_ ), .A2(_05425_ ), .ZN(_05426_ ) );
NAND2_X1 _12859_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][10] ), .ZN(_05427_ ) );
NAND2_X1 _12860_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][10] ), .ZN(_05428_ ) );
AOI21_X1 _12861_ ( .A(\fc_addr [15] ), .B1(_05427_ ), .B2(_05428_ ), .ZN(_05429_ ) );
AND3_X1 _12862_ ( .A1(_05427_ ), .A2(\fc_addr [15] ), .A3(_05428_ ), .ZN(_05430_ ) );
OR4_X1 _12863_ ( .A1(_05423_ ), .A2(_05426_ ), .A3(_05429_ ), .A4(_05430_ ), .ZN(_05431_ ) );
NAND2_X1 _12864_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][9] ), .ZN(_05432_ ) );
NAND2_X1 _12865_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][9] ), .ZN(_05433_ ) );
AOI21_X1 _12866_ ( .A(\fc_addr [14] ), .B1(_05432_ ), .B2(_05433_ ), .ZN(_05434_ ) );
AND3_X1 _12867_ ( .A1(_05432_ ), .A2(\fc_addr [14] ), .A3(_05433_ ), .ZN(_05435_ ) );
NAND2_X1 _12868_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][11] ), .ZN(_05436_ ) );
NAND2_X1 _12869_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][11] ), .ZN(_05437_ ) );
NAND2_X1 _12870_ ( .A1(_05436_ ), .A2(_05437_ ), .ZN(_05438_ ) );
INV_X1 _12871_ ( .A(\fc_addr [16] ), .ZN(_05439_ ) );
XNOR2_X1 _12872_ ( .A(_05438_ ), .B(_05439_ ), .ZN(_05440_ ) );
NOR4_X1 _12873_ ( .A1(_05431_ ), .A2(_05434_ ), .A3(_05435_ ), .A4(_05440_ ), .ZN(_05441_ ) );
INV_X1 _12874_ ( .A(\fc_addr [31] ), .ZN(_05442_ ) );
NAND2_X1 _12875_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][26] ), .ZN(_05443_ ) );
NAND2_X1 _12876_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][26] ), .ZN(_05444_ ) );
AOI21_X1 _12877_ ( .A(_05442_ ), .B1(_05443_ ), .B2(_05444_ ), .ZN(_05445_ ) );
AND3_X1 _12878_ ( .A1(_05443_ ), .A2(_05442_ ), .A3(_05444_ ), .ZN(_05446_ ) );
OAI211_X1 _12879_ ( .A(_05420_ ), .B(_05441_ ), .C1(_05445_ ), .C2(_05446_ ), .ZN(_05447_ ) );
MUX2_X1 _12880_ ( .A(\u_icache.ctags[0][16] ), .B(\u_icache.ctags[1][16] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05448_ ) );
XNOR2_X1 _12881_ ( .A(_05448_ ), .B(\fc_addr [21] ), .ZN(_05449_ ) );
MUX2_X1 _12882_ ( .A(\u_icache.ctags[0][17] ), .B(\u_icache.ctags[1][17] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05450_ ) );
INV_X1 _12883_ ( .A(\fc_addr [22] ), .ZN(_05451_ ) );
NAND2_X1 _12884_ ( .A1(_05450_ ), .A2(_05451_ ), .ZN(_05452_ ) );
NAND2_X1 _12885_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][19] ), .ZN(_05453_ ) );
NAND2_X1 _12886_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][19] ), .ZN(_05454_ ) );
NAND3_X1 _12887_ ( .A1(_05453_ ), .A2(\fc_addr [24] ), .A3(_05454_ ), .ZN(_05455_ ) );
AND3_X1 _12888_ ( .A1(_05449_ ), .A2(_05452_ ), .A3(_05455_ ), .ZN(_05456_ ) );
NAND2_X1 _12889_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][20] ), .ZN(_05457_ ) );
INV_X1 _12890_ ( .A(\fc_addr [25] ), .ZN(_05458_ ) );
NAND2_X1 _12891_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][20] ), .ZN(_05459_ ) );
AND3_X1 _12892_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(_05459_ ), .ZN(_05460_ ) );
AOI21_X1 _12893_ ( .A(_05458_ ), .B1(_05457_ ), .B2(_05459_ ), .ZN(_05461_ ) );
INV_X1 _12894_ ( .A(\fc_addr [27] ), .ZN(_05462_ ) );
NAND2_X1 _12895_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][22] ), .ZN(_05463_ ) );
NAND2_X1 _12896_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][22] ), .ZN(_05464_ ) );
AOI21_X1 _12897_ ( .A(_05462_ ), .B1(_05463_ ), .B2(_05464_ ), .ZN(_05465_ ) );
AND3_X1 _12898_ ( .A1(_05463_ ), .A2(_05462_ ), .A3(_05464_ ), .ZN(_05466_ ) );
OAI221_X1 _12899_ ( .A(_05456_ ), .B1(_05460_ ), .B2(_05461_ ), .C1(_05465_ ), .C2(_05466_ ), .ZN(_05467_ ) );
MUX2_X1 _12900_ ( .A(\u_icache.ctags[0][21] ), .B(\u_icache.ctags[1][21] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05468_ ) );
INV_X1 _12901_ ( .A(\fc_addr [26] ), .ZN(_05469_ ) );
AND2_X1 _12902_ ( .A1(_05468_ ), .A2(_05469_ ), .ZN(_05470_ ) );
NOR2_X1 _12903_ ( .A1(_05468_ ), .A2(_05469_ ), .ZN(_05471_ ) );
AND3_X1 _12904_ ( .A1(_05408_ ), .A2(\fc_addr [28] ), .A3(_05409_ ), .ZN(_05472_ ) );
AOI21_X1 _12905_ ( .A(\fc_addr [24] ), .B1(_05453_ ), .B2(_05454_ ), .ZN(_05473_ ) );
OR4_X1 _12906_ ( .A1(_05470_ ), .A2(_05471_ ), .A3(_05472_ ), .A4(_05473_ ), .ZN(_05474_ ) );
NAND2_X1 _12907_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][18] ), .ZN(_05475_ ) );
INV_X1 _12908_ ( .A(\fc_addr [23] ), .ZN(_05476_ ) );
NAND2_X1 _12909_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][18] ), .ZN(_05477_ ) );
AND3_X1 _12910_ ( .A1(_05475_ ), .A2(_05476_ ), .A3(_05477_ ), .ZN(_05478_ ) );
AOI21_X1 _12911_ ( .A(_05476_ ), .B1(_05475_ ), .B2(_05477_ ), .ZN(_05479_ ) );
OAI22_X1 _12912_ ( .A1(_05478_ ), .A2(_05479_ ), .B1(_05450_ ), .B2(_05451_ ), .ZN(_05480_ ) );
NOR4_X1 _12913_ ( .A1(_05447_ ), .A2(_05467_ ), .A3(_05474_ ), .A4(_05480_ ), .ZN(_05481_ ) );
OR2_X1 _12914_ ( .A1(_05424_ ), .A2(_05425_ ), .ZN(_05482_ ) );
INV_X1 _12915_ ( .A(\u_icache.cvalids [0] ), .ZN(_05483_ ) );
INV_X1 _12916_ ( .A(\u_icache.cvalids [1] ), .ZN(_05484_ ) );
MUX2_X1 _12917_ ( .A(_05483_ ), .B(_05484_ ), .S(fanout_net_8 ), .Z(_05485_ ) );
MUX2_X1 _12918_ ( .A(\u_icache.ctags[0][1] ), .B(\u_icache.ctags[1][1] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05486_ ) );
INV_X1 _12919_ ( .A(\fc_addr [6] ), .ZN(_05487_ ) );
AND2_X1 _12920_ ( .A1(_05486_ ), .A2(_05487_ ), .ZN(_05488_ ) );
NAND2_X1 _12921_ ( .A1(_05406_ ), .A2(\u_icache.ctags[0][0] ), .ZN(_05489_ ) );
NAND2_X1 _12922_ ( .A1(\u_icache.ctags[1][0] ), .A2(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .ZN(_05490_ ) );
AND3_X1 _12923_ ( .A1(_05489_ ), .A2(\fc_addr [5] ), .A3(_05490_ ), .ZN(_05491_ ) );
AOI21_X1 _12924_ ( .A(\fc_addr [5] ), .B1(_05489_ ), .B2(_05490_ ), .ZN(_05492_ ) );
OR4_X1 _12925_ ( .A1(_05485_ ), .A2(_05488_ ), .A3(_05491_ ), .A4(_05492_ ), .ZN(_05493_ ) );
NAND2_X1 _12926_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][3] ), .ZN(_05494_ ) );
NAND2_X1 _12927_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][3] ), .ZN(_05495_ ) );
NAND2_X1 _12928_ ( .A1(_05494_ ), .A2(_05495_ ), .ZN(_05496_ ) );
INV_X1 _12929_ ( .A(\fc_addr [8] ), .ZN(_05497_ ) );
XNOR2_X1 _12930_ ( .A(_05496_ ), .B(_05497_ ), .ZN(_05498_ ) );
NAND2_X1 _12931_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][2] ), .ZN(_05499_ ) );
NAND2_X1 _12932_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][2] ), .ZN(_05500_ ) );
AOI21_X1 _12933_ ( .A(\fc_addr [7] ), .B1(_05499_ ), .B2(_05500_ ), .ZN(_05501_ ) );
NOR2_X1 _12934_ ( .A1(_05486_ ), .A2(_05487_ ), .ZN(_05502_ ) );
NOR4_X1 _12935_ ( .A1(_05493_ ), .A2(_05498_ ), .A3(_05501_ ), .A4(_05502_ ), .ZN(_05503_ ) );
NAND2_X1 _12936_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][14] ), .ZN(_05504_ ) );
NAND2_X1 _12937_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][14] ), .ZN(_05505_ ) );
AND3_X1 _12938_ ( .A1(_05504_ ), .A2(\fc_addr [19] ), .A3(_05505_ ), .ZN(_05506_ ) );
NAND2_X1 _12939_ ( .A1(_05406_ ), .A2(\u_icache.ctags[0][4] ), .ZN(_05507_ ) );
NAND2_X1 _12940_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][4] ), .ZN(_05508_ ) );
AND3_X1 _12941_ ( .A1(_05507_ ), .A2(\fc_addr [9] ), .A3(_05508_ ), .ZN(_05509_ ) );
AOI21_X1 _12942_ ( .A(\fc_addr [17] ), .B1(_05421_ ), .B2(_05422_ ), .ZN(_05510_ ) );
AOI21_X1 _12943_ ( .A(\fc_addr [19] ), .B1(_05504_ ), .B2(_05505_ ), .ZN(_05511_ ) );
OR4_X1 _12944_ ( .A1(_05506_ ), .A2(_05509_ ), .A3(_05510_ ), .A4(_05511_ ), .ZN(_05512_ ) );
NAND2_X1 _12945_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][7] ), .ZN(_05513_ ) );
NAND2_X1 _12946_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][7] ), .ZN(_05514_ ) );
NAND2_X1 _12947_ ( .A1(_05513_ ), .A2(_05514_ ), .ZN(_05515_ ) );
INV_X1 _12948_ ( .A(\fc_addr [12] ), .ZN(_05516_ ) );
XNOR2_X1 _12949_ ( .A(_05515_ ), .B(_05516_ ), .ZN(_05517_ ) );
NAND2_X1 _12950_ ( .A1(_05407_ ), .A2(\u_icache.ctags[0][5] ), .ZN(_05518_ ) );
NAND2_X1 _12951_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][5] ), .ZN(_05519_ ) );
AOI21_X1 _12952_ ( .A(\fc_addr [10] ), .B1(_05518_ ), .B2(_05519_ ), .ZN(_05520_ ) );
AND3_X1 _12953_ ( .A1(_05518_ ), .A2(\fc_addr [10] ), .A3(_05519_ ), .ZN(_05521_ ) );
NOR4_X1 _12954_ ( .A1(_05512_ ), .A2(_05517_ ), .A3(_05520_ ), .A4(_05521_ ), .ZN(_05522_ ) );
AND2_X1 _12955_ ( .A1(_05503_ ), .A2(_05522_ ), .ZN(_05523_ ) );
NAND2_X1 _12956_ ( .A1(_05412_ ), .A2(_05413_ ), .ZN(_05524_ ) );
INV_X1 _12957_ ( .A(\fc_addr [30] ), .ZN(_05525_ ) );
NAND2_X1 _12958_ ( .A1(_05524_ ), .A2(_05525_ ), .ZN(_05526_ ) );
NAND2_X1 _12959_ ( .A1(_05411_ ), .A2(\u_icache.ctags[0][15] ), .ZN(_05527_ ) );
NAND2_X1 _12960_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[1][15] ), .ZN(_05528_ ) );
NAND2_X1 _12961_ ( .A1(_05527_ ), .A2(_05528_ ), .ZN(_05529_ ) );
INV_X1 _12962_ ( .A(\fc_addr [20] ), .ZN(_05530_ ) );
XNOR2_X1 _12963_ ( .A(_05529_ ), .B(_05530_ ), .ZN(_05531_ ) );
MUX2_X1 _12964_ ( .A(\u_icache.ctags[0][6] ), .B(\u_icache.ctags[1][6] ), .S(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .Z(_05532_ ) );
INV_X1 _12965_ ( .A(\fc_addr [11] ), .ZN(_05533_ ) );
NOR2_X1 _12966_ ( .A1(_05532_ ), .A2(_05533_ ), .ZN(_05534_ ) );
AND2_X1 _12967_ ( .A1(_05532_ ), .A2(_05533_ ), .ZN(_05535_ ) );
AOI21_X1 _12968_ ( .A(\fc_addr [9] ), .B1(_05507_ ), .B2(_05508_ ), .ZN(_05536_ ) );
AND3_X1 _12969_ ( .A1(_05499_ ), .A2(\fc_addr [7] ), .A3(_05500_ ), .ZN(_05537_ ) );
OR4_X1 _12970_ ( .A1(_05534_ ), .A2(_05535_ ), .A3(_05536_ ), .A4(_05537_ ), .ZN(_05538_ ) );
NOR2_X1 _12971_ ( .A1(_05411_ ), .A2(\u_icache.ctags[1][13] ), .ZN(_05539_ ) );
INV_X1 _12972_ ( .A(\fc_addr [18] ), .ZN(_05540_ ) );
NOR2_X1 _12973_ ( .A1(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .A2(\u_icache.ctags[0][13] ), .ZN(_05541_ ) );
OR3_X1 _12974_ ( .A1(_05539_ ), .A2(_05540_ ), .A3(_05541_ ), .ZN(_05542_ ) );
OAI21_X1 _12975_ ( .A(_05540_ ), .B1(_05539_ ), .B2(_05541_ ), .ZN(_05543_ ) );
AOI211_X1 _12976_ ( .A(_05531_ ), .B(_05538_ ), .C1(_05542_ ), .C2(_05543_ ), .ZN(_05544_ ) );
AND4_X1 _12977_ ( .A1(_05482_ ), .A2(_05523_ ), .A3(_05526_ ), .A4(_05544_ ), .ZN(_05545_ ) );
AOI211_X1 _12978_ ( .A(\u_icache.ended ), .B(_05405_ ), .C1(_05481_ ), .C2(_05545_ ), .ZN(_05546_ ) );
AND2_X1 _12979_ ( .A1(_05404_ ), .A2(_05546_ ), .ZN(_05547_ ) );
INV_X1 _12980_ ( .A(_00862_ ), .ZN(_05548_ ) );
NOR2_X1 _12981_ ( .A1(_05547_ ), .A2(_05548_ ), .ZN(_05549_ ) );
AND2_X1 _12982_ ( .A1(\u_lsu.rvalid ), .A2(\u_lsu.reading ), .ZN(_05550_ ) );
BUF_X2 _12983_ ( .A(_01145_ ), .Z(_05551_ ) );
AND2_X1 _12984_ ( .A1(_05550_ ), .A2(_05551_ ), .ZN(_05552_ ) );
AND2_X1 _12985_ ( .A1(_05549_ ), .A2(_05552_ ), .ZN(_05553_ ) );
AND3_X1 _12986_ ( .A1(\ca_addr [3] ), .A2(\ca_addr [4] ), .A3(\ca_addr [2] ), .ZN(_05554_ ) );
NAND3_X1 _12987_ ( .A1(_05554_ ), .A2(\ca_addr [5] ), .A3(\ca_addr [6] ), .ZN(_05555_ ) );
INV_X1 _12988_ ( .A(\ca_addr [7] ), .ZN(_05556_ ) );
NOR2_X1 _12989_ ( .A1(_05555_ ), .A2(_05556_ ), .ZN(_05557_ ) );
AND2_X1 _12990_ ( .A1(_05557_ ), .A2(\ca_addr [8] ), .ZN(_05558_ ) );
AND3_X1 _12991_ ( .A1(_05558_ ), .A2(\ca_addr [9] ), .A3(\ca_addr [10] ), .ZN(_05559_ ) );
AND2_X1 _12992_ ( .A1(_05559_ ), .A2(\ca_addr [11] ), .ZN(_05560_ ) );
AND2_X1 _12993_ ( .A1(_05560_ ), .A2(\ca_addr [12] ), .ZN(_05561_ ) );
AND3_X1 _12994_ ( .A1(_05561_ ), .A2(\ca_addr [14] ), .A3(\ca_addr [13] ), .ZN(_05562_ ) );
AND2_X1 _12995_ ( .A1(_05562_ ), .A2(\ca_addr [15] ), .ZN(_05563_ ) );
AND2_X1 _12996_ ( .A1(_05563_ ), .A2(\ca_addr [16] ), .ZN(_05564_ ) );
AND3_X1 _12997_ ( .A1(_05564_ ), .A2(\ca_addr [17] ), .A3(\ca_addr [18] ), .ZN(_05565_ ) );
AND2_X1 _12998_ ( .A1(_05565_ ), .A2(\ca_addr [19] ), .ZN(_05566_ ) );
AND2_X1 _12999_ ( .A1(_05566_ ), .A2(\ca_addr [20] ), .ZN(_05567_ ) );
AND2_X1 _13000_ ( .A1(\ca_addr [23] ), .A2(\ca_addr [22] ), .ZN(_05568_ ) );
AND4_X1 _13001_ ( .A1(\ca_addr [21] ), .A2(_05568_ ), .A3(\ca_addr [24] ), .A4(\ca_addr [25] ), .ZN(_05569_ ) );
NAND3_X1 _13002_ ( .A1(_05567_ ), .A2(\ca_addr [26] ), .A3(_05569_ ), .ZN(_05570_ ) );
INV_X1 _13003_ ( .A(\ca_addr [28] ), .ZN(_05571_ ) );
INV_X1 _13004_ ( .A(\ca_addr [27] ), .ZN(_05572_ ) );
NOR3_X1 _13005_ ( .A1(_05570_ ), .A2(_05571_ ), .A3(_05572_ ), .ZN(_05573_ ) );
AND3_X1 _13006_ ( .A1(_05573_ ), .A2(\ca_addr [29] ), .A3(\ca_addr [30] ), .ZN(_05574_ ) );
OAI21_X1 _13007_ ( .A(_05553_ ), .B1(_05574_ ), .B2(\ca_addr [31] ), .ZN(_05575_ ) );
AND4_X1 _13008_ ( .A1(\ca_addr [31] ), .A2(_05573_ ), .A3(\ca_addr [29] ), .A4(\ca_addr [30] ), .ZN(_05576_ ) );
AND2_X1 _13009_ ( .A1(_05547_ ), .A2(_00862_ ), .ZN(_00414_ ) );
INV_X2 _13010_ ( .A(_00414_ ), .ZN(_05577_ ) );
BUF_X4 _13011_ ( .A(_05577_ ), .Z(_05578_ ) );
OAI22_X1 _13012_ ( .A1(_05575_ ), .A2(_05576_ ), .B1(_05442_ ), .B2(_05578_ ), .ZN(_00336_ ) );
AOI22_X1 _13013_ ( .A1(_01100_ ), .A2(_01104_ ), .B1(_00758_ ), .B2(_01071_ ), .ZN(_05579_ ) );
AND2_X2 _13014_ ( .A1(_05579_ ), .A2(_01118_ ), .ZN(_05580_ ) );
NAND2_X1 _13015_ ( .A1(_01055_ ), .A2(_05580_ ), .ZN(_05581_ ) );
NOR3_X1 _13016_ ( .A1(_05581_ ), .A2(_00993_ ), .A3(_00916_ ), .ZN(_05582_ ) );
OAI21_X1 _13017_ ( .A(_05188_ ), .B1(_05582_ ), .B2(\u_exu.rlock [15] ), .ZN(_05583_ ) );
AND3_X1 _13018_ ( .A1(_01304_ ), .A2(_01289_ ), .A3(_01295_ ), .ZN(_05584_ ) );
AND3_X1 _13019_ ( .A1(_01286_ ), .A2(_01308_ ), .A3(_05584_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13020_ ( .A1(_05583_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00337_ ) );
BUF_X4 _13021_ ( .A(_04473_ ), .Z(_05585_ ) );
AND4_X1 _13022_ ( .A1(_01110_ ), .A2(_01107_ ), .A3(_00972_ ), .A4(_05580_ ), .ZN(_05586_ ) );
OAI21_X1 _13023_ ( .A(_05585_ ), .B1(_05586_ ), .B2(\u_exu.rlock [14] ), .ZN(_05587_ ) );
AND3_X1 _13024_ ( .A1(_01305_ ), .A2(_01289_ ), .A3(_01295_ ), .ZN(_05588_ ) );
AND3_X1 _13025_ ( .A1(_01286_ ), .A2(_01308_ ), .A3(_05588_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13026_ ( .A1(_05587_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ), .ZN(_00338_ ) );
NOR3_X1 _13027_ ( .A1(_05581_ ), .A2(_00920_ ), .A3(_00982_ ), .ZN(_05589_ ) );
OAI21_X1 _13028_ ( .A(_05585_ ), .B1(_05589_ ), .B2(\u_exu.rlock [5] ), .ZN(_05590_ ) );
BUF_X4 _13029_ ( .A(_01285_ ), .Z(_05591_ ) );
AND3_X1 _13030_ ( .A1(_01296_ ), .A2(_01304_ ), .A3(_01289_ ), .ZN(_05592_ ) );
INV_X1 _13031_ ( .A(_05592_ ), .ZN(_05593_ ) );
NOR3_X1 _13032_ ( .A1(_05591_ ), .A2(_01308_ ), .A3(_05593_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13033_ ( .A1(_05590_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00339_ ) );
NAND3_X1 _13034_ ( .A1(_01305_ ), .A2(_01296_ ), .A3(_01289_ ), .ZN(_05594_ ) );
NOR3_X1 _13035_ ( .A1(_05591_ ), .A2(_01308_ ), .A3(_05594_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_1_Y_$_AND__B_Y ) );
NAND4_X1 _13036_ ( .A1(_01107_ ), .A2(_01048_ ), .A3(_01110_ ), .A4(_05580_ ), .ZN(_05595_ ) );
AOI211_X1 _13037_ ( .A(_04460_ ), .B(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_1_Y_$_AND__B_Y ), .C1(_05595_ ), .C2(_01047_ ), .ZN(_00340_ ) );
AND4_X1 _13038_ ( .A1(_01110_ ), .A2(_01107_ ), .A3(_01009_ ), .A4(_05580_ ), .ZN(_05596_ ) );
OAI21_X1 _13039_ ( .A(_05585_ ), .B1(_05596_ ), .B2(\u_exu.rlock [3] ), .ZN(_05597_ ) );
AND3_X1 _13040_ ( .A1(_01290_ ), .A2(_01304_ ), .A3(_01295_ ), .ZN(_05598_ ) );
INV_X1 _13041_ ( .A(_05598_ ), .ZN(_05599_ ) );
NOR3_X1 _13042_ ( .A1(_05591_ ), .A2(_01308_ ), .A3(_05599_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13043_ ( .A1(_05597_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .ZN(_00341_ ) );
AND4_X1 _13044_ ( .A1(_01031_ ), .A2(_01107_ ), .A3(_01110_ ), .A4(_05580_ ), .ZN(_05600_ ) );
OAI21_X1 _13045_ ( .A(_05585_ ), .B1(_05600_ ), .B2(\u_exu.rlock [2] ), .ZN(_05601_ ) );
NOR3_X1 _13046_ ( .A1(_01296_ ), .A2(_01304_ ), .A3(_01289_ ), .ZN(_05602_ ) );
INV_X1 _13047_ ( .A(_05602_ ), .ZN(_05603_ ) );
NOR3_X1 _13048_ ( .A1(_05591_ ), .A2(_01308_ ), .A3(_05603_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13049_ ( .A1(_05601_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_00342_ ) );
NOR3_X1 _13050_ ( .A1(_05581_ ), .A2(_00920_ ), .A3(_00992_ ), .ZN(_05604_ ) );
OAI21_X1 _13051_ ( .A(_05585_ ), .B1(_05604_ ), .B2(\u_exu.rlock [1] ), .ZN(_05605_ ) );
NOR3_X1 _13052_ ( .A1(_01305_ ), .A2(_01289_ ), .A3(_01295_ ), .ZN(_05606_ ) );
INV_X1 _13053_ ( .A(_05606_ ), .ZN(_05607_ ) );
NOR3_X1 _13054_ ( .A1(_05591_ ), .A2(_01308_ ), .A3(_05607_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13055_ ( .A1(_05605_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .ZN(_00343_ ) );
AND4_X4 _13056_ ( .A1(_03740_ ), .A2(_03739_ ), .A3(_00985_ ), .A4(_05580_ ), .ZN(_05608_ ) );
OAI21_X1 _13057_ ( .A(_04476_ ), .B1(_05608_ ), .B2(\u_exu.rlock [0] ), .ZN(_05609_ ) );
NOR3_X1 _13058_ ( .A1(_01304_ ), .A2(_01289_ ), .A3(_01295_ ), .ZN(_05610_ ) );
AND2_X1 _13059_ ( .A1(_05610_ ), .A2(_01300_ ), .ZN(_05611_ ) );
AOI21_X1 _13060_ ( .A(_05609_ ), .B1(_01286_ ), .B2(_05611_ ), .ZN(_00344_ ) );
AND4_X1 _13061_ ( .A1(_01110_ ), .A2(_01107_ ), .A3(_00999_ ), .A4(_05580_ ), .ZN(_05612_ ) );
OAI21_X1 _13062_ ( .A(_05585_ ), .B1(_05612_ ), .B2(\u_exu.rlock [13] ), .ZN(_05613_ ) );
NOR3_X1 _13063_ ( .A1(_05591_ ), .A2(_01300_ ), .A3(_05593_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13064_ ( .A1(_05613_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_00345_ ) );
NOR3_X1 _13065_ ( .A1(_05581_ ), .A2(_00993_ ), .A3(_01021_ ), .ZN(_05614_ ) );
OAI21_X1 _13066_ ( .A(_05585_ ), .B1(_05614_ ), .B2(\u_exu.rlock [12] ), .ZN(_05615_ ) );
NOR3_X1 _13067_ ( .A1(_05591_ ), .A2(_01300_ ), .A3(_05594_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13068_ ( .A1(_05615_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ), .ZN(_00346_ ) );
NOR3_X1 _13069_ ( .A1(_05581_ ), .A2(_00993_ ), .A3(_01008_ ), .ZN(_05616_ ) );
OAI21_X1 _13070_ ( .A(_05585_ ), .B1(_05616_ ), .B2(\u_exu.rlock [11] ), .ZN(_05617_ ) );
NOR3_X1 _13071_ ( .A1(_05591_ ), .A2(_01300_ ), .A3(_05599_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13072_ ( .A1(_05617_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_00347_ ) );
NOR3_X1 _13073_ ( .A1(_05581_ ), .A2(_00993_ ), .A3(_01013_ ), .ZN(_05618_ ) );
OAI21_X1 _13074_ ( .A(_05585_ ), .B1(_05618_ ), .B2(\u_exu.rlock [10] ), .ZN(_05619_ ) );
NOR3_X1 _13075_ ( .A1(_05591_ ), .A2(_01300_ ), .A3(_05603_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13076_ ( .A1(_05619_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_00348_ ) );
AND4_X1 _13077_ ( .A1(_01110_ ), .A2(_01107_ ), .A3(_00994_ ), .A4(_05580_ ), .ZN(_05620_ ) );
OAI21_X1 _13078_ ( .A(_05585_ ), .B1(_05620_ ), .B2(\u_exu.rlock [9] ), .ZN(_05621_ ) );
NOR3_X1 _13079_ ( .A1(_05591_ ), .A2(_01300_ ), .A3(_05607_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13080_ ( .A1(_05621_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_00349_ ) );
BUF_X4 _13081_ ( .A(_04473_ ), .Z(_05622_ ) );
AND4_X1 _13082_ ( .A1(_01110_ ), .A2(_01107_ ), .A3(_00963_ ), .A4(_05580_ ), .ZN(_05623_ ) );
OAI21_X1 _13083_ ( .A(_05622_ ), .B1(_05623_ ), .B2(\u_exu.rlock [8] ), .ZN(_05624_ ) );
AND3_X1 _13084_ ( .A1(_01286_ ), .A2(_01308_ ), .A3(_05610_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13085_ ( .A1(_05624_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ), .ZN(_00350_ ) );
NOR3_X1 _13086_ ( .A1(_05581_ ), .A2(_00920_ ), .A3(_00916_ ), .ZN(_05625_ ) );
OAI21_X1 _13087_ ( .A(_05622_ ), .B1(_05625_ ), .B2(\u_exu.rlock [7] ), .ZN(_05626_ ) );
AND3_X1 _13088_ ( .A1(_01286_ ), .A2(_01300_ ), .A3(_05584_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13089_ ( .A1(_05626_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_00351_ ) );
AND4_X1 _13090_ ( .A1(_01036_ ), .A2(_01107_ ), .A3(_01110_ ), .A4(_05580_ ), .ZN(_05627_ ) );
OAI21_X1 _13091_ ( .A(_05622_ ), .B1(_05627_ ), .B2(\u_exu.rlock [6] ), .ZN(_05628_ ) );
AND3_X1 _13092_ ( .A1(_01286_ ), .A2(_01300_ ), .A3(_05588_ ), .ZN(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _13093_ ( .A1(_05628_ ), .A2(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00352_ ) );
INV_X1 _13094_ ( .A(_05553_ ), .ZN(_05629_ ) );
BUF_X4 _13095_ ( .A(_05629_ ), .Z(_05630_ ) );
NAND4_X1 _13096_ ( .A1(\ca_addr [23] ), .A2(\ca_addr [22] ), .A3(\ca_addr [21] ), .A4(\ca_addr [25] ), .ZN(_05631_ ) );
INV_X1 _13097_ ( .A(\ca_addr [24] ), .ZN(_05632_ ) );
INV_X1 _13098_ ( .A(\ca_addr [20] ), .ZN(_05633_ ) );
NOR3_X1 _13099_ ( .A1(_05631_ ), .A2(_05632_ ), .A3(_05633_ ), .ZN(_05634_ ) );
NAND3_X1 _13100_ ( .A1(_05566_ ), .A2(\ca_addr [26] ), .A3(_05634_ ), .ZN(_05635_ ) );
NOR2_X1 _13101_ ( .A1(_05635_ ), .A2(_05572_ ), .ZN(_05636_ ) );
AND3_X1 _13102_ ( .A1(_05636_ ), .A2(\ca_addr [29] ), .A3(\ca_addr [28] ), .ZN(_05637_ ) );
XNOR2_X1 _13103_ ( .A(_05637_ ), .B(\ca_addr [30] ), .ZN(_05638_ ) );
OAI22_X1 _13104_ ( .A1(_05630_ ), .A2(_05638_ ), .B1(_05525_ ), .B2(_05578_ ), .ZN(_00353_ ) );
BUF_X4 _13105_ ( .A(_05549_ ), .Z(_05639_ ) );
BUF_X4 _13106_ ( .A(_05552_ ), .Z(_05640_ ) );
BUF_X2 _13107_ ( .A(_05640_ ), .Z(icah_ready ) );
AND2_X1 _13108_ ( .A1(_05558_ ), .A2(\ca_addr [9] ), .ZN(_05641_ ) );
AND4_X1 _13109_ ( .A1(\ca_addr [16] ), .A2(\ca_addr [14] ), .A3(\ca_addr [15] ), .A4(\ca_addr [17] ), .ZN(_05642_ ) );
AND2_X1 _13110_ ( .A1(\ca_addr [11] ), .A2(\ca_addr [10] ), .ZN(_05643_ ) );
AND4_X1 _13111_ ( .A1(\ca_addr [13] ), .A2(_05642_ ), .A3(\ca_addr [12] ), .A4(_05643_ ), .ZN(_05644_ ) );
AND2_X1 _13112_ ( .A1(_05641_ ), .A2(_05644_ ), .ZN(_05645_ ) );
AND3_X1 _13113_ ( .A1(_05645_ ), .A2(\ca_addr [19] ), .A3(\ca_addr [18] ), .ZN(_05646_ ) );
AND2_X1 _13114_ ( .A1(_05646_ ), .A2(\ca_addr [20] ), .ZN(_05647_ ) );
OAI211_X1 _13115_ ( .A(_05639_ ), .B(icah_ready ), .C1(\ca_addr [21] ), .C2(_05647_ ), .ZN(_05648_ ) );
AND2_X1 _13116_ ( .A1(_05567_ ), .A2(\ca_addr [21] ), .ZN(_05649_ ) );
INV_X1 _13117_ ( .A(\fc_addr [21] ), .ZN(_05650_ ) );
OAI22_X1 _13118_ ( .A1(_05648_ ), .A2(_05649_ ), .B1(_05650_ ), .B2(_05578_ ), .ZN(_00354_ ) );
OAI211_X1 _13119_ ( .A(_05639_ ), .B(icah_ready ), .C1(\ca_addr [20] ), .C2(_05646_ ), .ZN(_05651_ ) );
OAI22_X1 _13120_ ( .A1(_05651_ ), .A2(_05567_ ), .B1(_05530_ ), .B2(_05578_ ), .ZN(_00355_ ) );
AND4_X1 _13121_ ( .A1(\ca_addr [9] ), .A2(_05558_ ), .A3(\ca_addr [18] ), .A4(_05644_ ), .ZN(_05652_ ) );
OAI211_X1 _13122_ ( .A(_05639_ ), .B(icah_ready ), .C1(\ca_addr [19] ), .C2(_05652_ ), .ZN(_05653_ ) );
INV_X1 _13123_ ( .A(\fc_addr [19] ), .ZN(_05654_ ) );
OAI22_X1 _13124_ ( .A1(_05653_ ), .A2(_05566_ ), .B1(_05654_ ), .B2(_05578_ ), .ZN(_00356_ ) );
XOR2_X1 _13125_ ( .A(_05645_ ), .B(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_B ), .Z(_05655_ ) );
OAI22_X1 _13126_ ( .A1(_05630_ ), .A2(_05655_ ), .B1(_05540_ ), .B2(_05578_ ), .ZN(_00357_ ) );
XNOR2_X1 _13127_ ( .A(_05564_ ), .B(\ca_addr [17] ), .ZN(_05656_ ) );
INV_X1 _13128_ ( .A(\fc_addr [17] ), .ZN(_05657_ ) );
BUF_X4 _13129_ ( .A(_05577_ ), .Z(_05658_ ) );
OAI22_X1 _13130_ ( .A1(_05630_ ), .A2(_05656_ ), .B1(_05657_ ), .B2(_05658_ ), .ZN(_00358_ ) );
OAI211_X1 _13131_ ( .A(_05639_ ), .B(icah_ready ), .C1(\ca_addr [16] ), .C2(_05563_ ), .ZN(_05659_ ) );
OAI22_X1 _13132_ ( .A1(_05659_ ), .A2(_05564_ ), .B1(_05439_ ), .B2(_05658_ ), .ZN(_00359_ ) );
XNOR2_X1 _13133_ ( .A(_05562_ ), .B(\ca_addr [15] ), .ZN(_05660_ ) );
INV_X1 _13134_ ( .A(\fc_addr [15] ), .ZN(_05661_ ) );
OAI22_X1 _13135_ ( .A1(_05630_ ), .A2(_05660_ ), .B1(_05661_ ), .B2(_05658_ ), .ZN(_00360_ ) );
AND2_X1 _13136_ ( .A1(_05561_ ), .A2(\ca_addr [13] ), .ZN(_05662_ ) );
XNOR2_X1 _13137_ ( .A(_05662_ ), .B(\ca_addr [14] ), .ZN(_05663_ ) );
INV_X1 _13138_ ( .A(\fc_addr [14] ), .ZN(_05664_ ) );
OAI22_X1 _13139_ ( .A1(_05630_ ), .A2(_05663_ ), .B1(_05664_ ), .B2(_05658_ ), .ZN(_00361_ ) );
AND3_X1 _13140_ ( .A1(_05641_ ), .A2(\ca_addr [12] ), .A3(_05643_ ), .ZN(_05665_ ) );
OAI211_X1 _13141_ ( .A(_05639_ ), .B(icah_ready ), .C1(\ca_addr [13] ), .C2(_05665_ ), .ZN(_05666_ ) );
OAI22_X1 _13142_ ( .A1(_05666_ ), .A2(_05662_ ), .B1(_05425_ ), .B2(_05658_ ), .ZN(_00362_ ) );
OAI211_X1 _13143_ ( .A(_05639_ ), .B(icah_ready ), .C1(\ca_addr [12] ), .C2(_05560_ ), .ZN(_05667_ ) );
OAI22_X1 _13144_ ( .A1(_05667_ ), .A2(_05561_ ), .B1(_05516_ ), .B2(_05658_ ), .ZN(_00363_ ) );
AND4_X1 _13145_ ( .A1(\ca_addr [19] ), .A2(\ca_addr [21] ), .A3(\ca_addr [20] ), .A4(\ca_addr [18] ), .ZN(_05668_ ) );
AND4_X1 _13146_ ( .A1(\ca_addr [24] ), .A2(_05668_ ), .A3(\ca_addr [25] ), .A4(_05568_ ), .ZN(_05669_ ) );
AND2_X1 _13147_ ( .A1(_05645_ ), .A2(_05669_ ), .ZN(_05670_ ) );
NAND3_X1 _13148_ ( .A1(_05670_ ), .A2(\ca_addr [27] ), .A3(\ca_addr [26] ), .ZN(_05671_ ) );
NOR2_X1 _13149_ ( .A1(_05671_ ), .A2(_05571_ ), .ZN(_05672_ ) );
OAI211_X1 _13150_ ( .A(_05639_ ), .B(_05640_ ), .C1(\ca_addr [29] ), .C2(_05672_ ), .ZN(_05673_ ) );
OAI22_X1 _13151_ ( .A1(_05673_ ), .A2(_05637_ ), .B1(_05416_ ), .B2(_05658_ ), .ZN(_00364_ ) );
XNOR2_X1 _13152_ ( .A(_05559_ ), .B(\ca_addr [11] ), .ZN(_05674_ ) );
OAI22_X1 _13153_ ( .A1(_05630_ ), .A2(_05674_ ), .B1(_05533_ ), .B2(_05658_ ), .ZN(_00365_ ) );
XOR2_X1 _13154_ ( .A(_05641_ ), .B(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_B ), .Z(_05675_ ) );
INV_X1 _13155_ ( .A(\fc_addr [10] ), .ZN(_05676_ ) );
OAI22_X1 _13156_ ( .A1(_05630_ ), .A2(_05675_ ), .B1(_05676_ ), .B2(_05658_ ), .ZN(_00366_ ) );
XNOR2_X1 _13157_ ( .A(_05558_ ), .B(\ca_addr [9] ), .ZN(_05677_ ) );
INV_X1 _13158_ ( .A(\fc_addr [9] ), .ZN(_05678_ ) );
OAI22_X1 _13159_ ( .A1(_05630_ ), .A2(_05677_ ), .B1(_05678_ ), .B2(_05658_ ), .ZN(_00367_ ) );
XOR2_X1 _13160_ ( .A(_05557_ ), .B(\u_icache.caddr_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ), .Z(_05679_ ) );
OAI22_X1 _13161_ ( .A1(_05630_ ), .A2(_05679_ ), .B1(_05497_ ), .B2(_05577_ ), .ZN(_00368_ ) );
XNOR2_X1 _13162_ ( .A(_05555_ ), .B(_05556_ ), .ZN(_05680_ ) );
INV_X1 _13163_ ( .A(\fc_addr [7] ), .ZN(_05681_ ) );
OAI22_X1 _13164_ ( .A1(_05630_ ), .A2(_05680_ ), .B1(_05681_ ), .B2(_05577_ ), .ZN(_00369_ ) );
AND2_X1 _13165_ ( .A1(_05554_ ), .A2(\ca_addr [5] ), .ZN(_05682_ ) );
XOR2_X1 _13166_ ( .A(_05682_ ), .B(\u_icache.caddr_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ), .Z(_05683_ ) );
OAI22_X1 _13167_ ( .A1(_05629_ ), .A2(_05683_ ), .B1(_05487_ ), .B2(_05577_ ), .ZN(_00370_ ) );
OAI211_X1 _13168_ ( .A(_05639_ ), .B(_05640_ ), .C1(\ca_addr [5] ), .C2(_05554_ ), .ZN(_05684_ ) );
INV_X1 _13169_ ( .A(\fc_addr [5] ), .ZN(_05685_ ) );
OAI22_X1 _13170_ ( .A1(_05684_ ), .A2(_05682_ ), .B1(_05685_ ), .B2(_05577_ ), .ZN(_00371_ ) );
AND2_X1 _13171_ ( .A1(\ca_addr [3] ), .A2(\ca_addr [2] ), .ZN(_05686_ ) );
XOR2_X1 _13172_ ( .A(_05686_ ), .B(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_B ), .Z(_05687_ ) );
INV_X4 _13173_ ( .A(fanout_net_8 ), .ZN(_05688_ ) );
BUF_X4 _13174_ ( .A(_05688_ ), .Z(_05689_ ) );
BUF_X4 _13175_ ( .A(_05689_ ), .Z(_05690_ ) );
OAI22_X1 _13176_ ( .A1(_05629_ ), .A2(_05687_ ), .B1(_05690_ ), .B2(_05577_ ), .ZN(_00372_ ) );
NOR2_X1 _13177_ ( .A1(\ca_addr [3] ), .A2(\ca_addr [2] ), .ZN(_05691_ ) );
NOR4_X1 _13178_ ( .A1(_05547_ ), .A2(_05548_ ), .A3(_05686_ ), .A4(_05691_ ), .ZN(_00373_ ) );
AOI211_X1 _13179_ ( .A(_01210_ ), .B(_05548_ ), .C1(_05404_ ), .C2(_05546_ ), .ZN(_00374_ ) );
XNOR2_X1 _13180_ ( .A(_05671_ ), .B(_05571_ ), .ZN(_05692_ ) );
INV_X1 _13181_ ( .A(\fc_addr [28] ), .ZN(_05693_ ) );
OAI22_X1 _13182_ ( .A1(_05629_ ), .A2(_05692_ ), .B1(_05693_ ), .B2(_05577_ ), .ZN(_00375_ ) );
AND4_X1 _13183_ ( .A1(\ca_addr [26] ), .A2(_05641_ ), .A3(_05644_ ), .A4(_05669_ ), .ZN(_05694_ ) );
OAI211_X1 _13184_ ( .A(_05639_ ), .B(_05640_ ), .C1(\ca_addr [27] ), .C2(_05694_ ), .ZN(_05695_ ) );
OAI22_X1 _13185_ ( .A1(_05695_ ), .A2(_05636_ ), .B1(_05462_ ), .B2(_05577_ ), .ZN(_00376_ ) );
OAI211_X1 _13186_ ( .A(_05639_ ), .B(_05640_ ), .C1(_01178_ ), .C2(_05670_ ), .ZN(_05696_ ) );
AND4_X1 _13187_ ( .A1(\ca_addr [20] ), .A2(_05566_ ), .A3(_01178_ ), .A4(_05569_ ), .ZN(_05697_ ) );
OAI22_X1 _13188_ ( .A1(_05696_ ), .A2(_05697_ ), .B1(_05469_ ), .B2(_05577_ ), .ZN(_00377_ ) );
INV_X1 _13189_ ( .A(_05547_ ), .ZN(_05698_ ) );
AND2_X1 _13190_ ( .A1(_05567_ ), .A2(_05569_ ), .ZN(_05699_ ) );
INV_X1 _13191_ ( .A(_05699_ ), .ZN(_05700_ ) );
NAND4_X1 _13192_ ( .A1(_05698_ ), .A2(_00863_ ), .A3(_05700_ ), .A4(_05640_ ), .ZN(_05701_ ) );
AND3_X1 _13193_ ( .A1(_05647_ ), .A2(\ca_addr [21] ), .A3(_05568_ ), .ZN(_05702_ ) );
AOI21_X1 _13194_ ( .A(\ca_addr [25] ), .B1(_05702_ ), .B2(\ca_addr [24] ), .ZN(_05703_ ) );
OAI22_X1 _13195_ ( .A1(_05578_ ), .A2(_05458_ ), .B1(_05701_ ), .B2(_05703_ ), .ZN(_00378_ ) );
AND3_X1 _13196_ ( .A1(_05567_ ), .A2(\ca_addr [21] ), .A3(_05568_ ), .ZN(_05704_ ) );
NAND2_X1 _13197_ ( .A1(_05704_ ), .A2(\ca_addr [24] ), .ZN(_05705_ ) );
NAND4_X1 _13198_ ( .A1(_05705_ ), .A2(_05698_ ), .A3(_05640_ ), .A4(_00863_ ), .ZN(_05706_ ) );
NOR2_X1 _13199_ ( .A1(_05702_ ), .A2(\ca_addr [24] ), .ZN(_05707_ ) );
INV_X1 _13200_ ( .A(\fc_addr [24] ), .ZN(_05708_ ) );
OAI22_X1 _13201_ ( .A1(_05706_ ), .A2(_05707_ ), .B1(_05578_ ), .B2(_05708_ ), .ZN(_00379_ ) );
INV_X1 _13202_ ( .A(_05704_ ), .ZN(_05709_ ) );
NAND4_X1 _13203_ ( .A1(_05698_ ), .A2(_05709_ ), .A3(_00863_ ), .A4(_05640_ ), .ZN(_05710_ ) );
AND3_X1 _13204_ ( .A1(_05647_ ), .A2(\ca_addr [22] ), .A3(\ca_addr [21] ), .ZN(_05711_ ) );
NOR2_X1 _13205_ ( .A1(_05711_ ), .A2(\ca_addr [23] ), .ZN(_05712_ ) );
OAI22_X1 _13206_ ( .A1(_05710_ ), .A2(_05712_ ), .B1(_05578_ ), .B2(_05476_ ), .ZN(_00380_ ) );
AND3_X1 _13207_ ( .A1(_05567_ ), .A2(\ca_addr [22] ), .A3(\ca_addr [21] ), .ZN(_05713_ ) );
INV_X1 _13208_ ( .A(_05713_ ), .ZN(_05714_ ) );
NAND4_X1 _13209_ ( .A1(_05698_ ), .A2(_05714_ ), .A3(_05640_ ), .A4(_00863_ ), .ZN(_05715_ ) );
AOI21_X1 _13210_ ( .A(\ca_addr [22] ), .B1(_05647_ ), .B2(\ca_addr [21] ), .ZN(_05716_ ) );
OAI22_X1 _13211_ ( .A1(_05715_ ), .A2(_05716_ ), .B1(_05578_ ), .B2(_05451_ ), .ZN(_00381_ ) );
BUF_X4 _13212_ ( .A(_00764_ ), .Z(_05717_ ) );
BUF_X4 _13213_ ( .A(_05717_ ), .Z(_05718_ ) );
INV_X1 _13214_ ( .A(fanout_net_6 ), .ZN(_05719_ ) );
CLKBUF_X2 _13215_ ( .A(_05719_ ), .Z(_05720_ ) );
CLKBUF_X3 _13216_ ( .A(_05720_ ), .Z(_05721_ ) );
OR2_X1 _13217_ ( .A1(_05721_ ), .A2(\u_icache.cblocks[1][31] ), .ZN(_05722_ ) );
INV_X1 _13218_ ( .A(\fc_addr [3] ), .ZN(_05723_ ) );
BUF_X4 _13219_ ( .A(_05723_ ), .Z(_05724_ ) );
BUF_X4 _13220_ ( .A(_05724_ ), .Z(_05725_ ) );
OAI211_X1 _13221_ ( .A(_05722_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][31] ), .ZN(_05726_ ) );
NOR2_X2 _13222_ ( .A1(_05723_ ), .A2(fanout_net_6 ), .ZN(_05727_ ) );
BUF_X4 _13223_ ( .A(_05727_ ), .Z(_05728_ ) );
AND2_X2 _13224_ ( .A1(\fc_addr [3] ), .A2(fanout_net_6 ), .ZN(_05729_ ) );
BUF_X4 _13225_ ( .A(_05729_ ), .Z(_05730_ ) );
BUF_X4 _13226_ ( .A(_05730_ ), .Z(_05731_ ) );
AOI22_X1 _13227_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][31] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][31] ), .ZN(_05732_ ) );
AOI21_X1 _13228_ ( .A(fanout_net_8 ), .B1(_05726_ ), .B2(_05732_ ), .ZN(_05733_ ) );
CLKBUF_X2 _13229_ ( .A(_05720_ ), .Z(_05734_ ) );
OR2_X1 _13230_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[5][31] ), .ZN(_05735_ ) );
BUF_X4 _13231_ ( .A(_05724_ ), .Z(_05736_ ) );
OAI211_X1 _13232_ ( .A(_05735_ ), .B(_05736_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][31] ), .ZN(_05737_ ) );
BUF_X4 _13233_ ( .A(_05727_ ), .Z(_05738_ ) );
BUF_X4 _13234_ ( .A(_05730_ ), .Z(_05739_ ) );
AOI22_X1 _13235_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[6][31] ), .B1(_05739_ ), .B2(\u_icache.cblocks[7][31] ), .ZN(_05740_ ) );
AOI21_X1 _13236_ ( .A(_05690_ ), .B1(_05737_ ), .B2(_05740_ ), .ZN(_05741_ ) );
NOR2_X1 _13237_ ( .A1(_05733_ ), .A2(_05741_ ), .ZN(_05742_ ) );
NOR3_X1 _13238_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05742_ ), .ZN(_00382_ ) );
OR2_X1 _13239_ ( .A1(_05721_ ), .A2(\u_icache.cblocks[1][30] ), .ZN(_05743_ ) );
OAI211_X1 _13240_ ( .A(_05743_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][30] ), .ZN(_05744_ ) );
AOI22_X1 _13241_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][30] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][30] ), .ZN(_05745_ ) );
AOI21_X1 _13242_ ( .A(fanout_net_8 ), .B1(_05744_ ), .B2(_05745_ ), .ZN(_05746_ ) );
BUF_X4 _13243_ ( .A(_05689_ ), .Z(_05747_ ) );
OR2_X1 _13244_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[5][30] ), .ZN(_05748_ ) );
OAI211_X1 _13245_ ( .A(_05748_ ), .B(_05736_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][30] ), .ZN(_05749_ ) );
AOI22_X1 _13246_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[6][30] ), .B1(_05739_ ), .B2(\u_icache.cblocks[7][30] ), .ZN(_05750_ ) );
AOI21_X1 _13247_ ( .A(_05747_ ), .B1(_05749_ ), .B2(_05750_ ), .ZN(_05751_ ) );
NOR2_X1 _13248_ ( .A1(_05746_ ), .A2(_05751_ ), .ZN(_05752_ ) );
NOR3_X1 _13249_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05752_ ), .ZN(_00383_ ) );
OR2_X1 _13250_ ( .A1(_05721_ ), .A2(\u_icache.cblocks[1][21] ), .ZN(_05753_ ) );
OAI211_X1 _13251_ ( .A(_05753_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][21] ), .ZN(_05754_ ) );
AOI22_X1 _13252_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][21] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][21] ), .ZN(_05755_ ) );
AOI21_X1 _13253_ ( .A(fanout_net_8 ), .B1(_05754_ ), .B2(_05755_ ), .ZN(_05756_ ) );
OR2_X1 _13254_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[5][21] ), .ZN(_05757_ ) );
OAI211_X1 _13255_ ( .A(_05757_ ), .B(_05736_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][21] ), .ZN(_05758_ ) );
AOI22_X1 _13256_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[6][21] ), .B1(_05739_ ), .B2(\u_icache.cblocks[7][21] ), .ZN(_05759_ ) );
AOI21_X1 _13257_ ( .A(_05747_ ), .B1(_05758_ ), .B2(_05759_ ), .ZN(_05760_ ) );
NOR2_X1 _13258_ ( .A1(_05756_ ), .A2(_05760_ ), .ZN(_05761_ ) );
NOR3_X1 _13259_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05761_ ), .ZN(_00384_ ) );
OR2_X1 _13260_ ( .A1(_05721_ ), .A2(\u_icache.cblocks[1][20] ), .ZN(_05762_ ) );
OAI211_X1 _13261_ ( .A(_05762_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][20] ), .ZN(_05763_ ) );
AOI22_X1 _13262_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][20] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][20] ), .ZN(_05764_ ) );
AOI21_X1 _13263_ ( .A(fanout_net_8 ), .B1(_05763_ ), .B2(_05764_ ), .ZN(_05765_ ) );
CLKBUF_X2 _13264_ ( .A(_05720_ ), .Z(_05766_ ) );
OR2_X1 _13265_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][20] ), .ZN(_05767_ ) );
OAI211_X1 _13266_ ( .A(_05767_ ), .B(_05736_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][20] ), .ZN(_05768_ ) );
BUF_X4 _13267_ ( .A(_05730_ ), .Z(_05769_ ) );
AOI22_X1 _13268_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[6][20] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][20] ), .ZN(_05770_ ) );
AOI21_X1 _13269_ ( .A(_05747_ ), .B1(_05768_ ), .B2(_05770_ ), .ZN(_05771_ ) );
NOR2_X1 _13270_ ( .A1(_05765_ ), .A2(_05771_ ), .ZN(_05772_ ) );
NOR3_X1 _13271_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05772_ ), .ZN(_00385_ ) );
OR2_X1 _13272_ ( .A1(_05721_ ), .A2(\u_icache.cblocks[1][19] ), .ZN(_05773_ ) );
OAI211_X1 _13273_ ( .A(_05773_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][19] ), .ZN(_05774_ ) );
AOI22_X1 _13274_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][19] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][19] ), .ZN(_05775_ ) );
AOI21_X1 _13275_ ( .A(fanout_net_8 ), .B1(_05774_ ), .B2(_05775_ ), .ZN(_05776_ ) );
OR2_X1 _13276_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][19] ), .ZN(_05777_ ) );
OAI211_X1 _13277_ ( .A(_05777_ ), .B(_05736_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][19] ), .ZN(_05778_ ) );
BUF_X4 _13278_ ( .A(_05727_ ), .Z(_05779_ ) );
AOI22_X1 _13279_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][19] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][19] ), .ZN(_05780_ ) );
AOI21_X1 _13280_ ( .A(_05747_ ), .B1(_05778_ ), .B2(_05780_ ), .ZN(_05781_ ) );
NOR2_X1 _13281_ ( .A1(_05776_ ), .A2(_05781_ ), .ZN(_05782_ ) );
NOR3_X1 _13282_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05782_ ), .ZN(_00386_ ) );
CLKBUF_X2 _13283_ ( .A(_05720_ ), .Z(_05783_ ) );
OR2_X1 _13284_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][18] ), .ZN(_05784_ ) );
OAI211_X1 _13285_ ( .A(_05784_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][18] ), .ZN(_05785_ ) );
AOI22_X1 _13286_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][18] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][18] ), .ZN(_05786_ ) );
AOI21_X1 _13287_ ( .A(fanout_net_8 ), .B1(_05785_ ), .B2(_05786_ ), .ZN(_05787_ ) );
OR2_X1 _13288_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][18] ), .ZN(_05788_ ) );
OAI211_X1 _13289_ ( .A(_05788_ ), .B(_05736_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][18] ), .ZN(_05789_ ) );
AOI22_X1 _13290_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][18] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][18] ), .ZN(_05790_ ) );
AOI21_X1 _13291_ ( .A(_05747_ ), .B1(_05789_ ), .B2(_05790_ ), .ZN(_05791_ ) );
NOR2_X1 _13292_ ( .A1(_05787_ ), .A2(_05791_ ), .ZN(_05792_ ) );
NOR3_X1 _13293_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05792_ ), .ZN(_00387_ ) );
OR2_X1 _13294_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][17] ), .ZN(_05793_ ) );
OAI211_X1 _13295_ ( .A(_05793_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][17] ), .ZN(_05794_ ) );
AOI22_X1 _13296_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][17] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][17] ), .ZN(_05795_ ) );
AOI21_X1 _13297_ ( .A(fanout_net_8 ), .B1(_05794_ ), .B2(_05795_ ), .ZN(_05796_ ) );
OR2_X1 _13298_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][17] ), .ZN(_05797_ ) );
OAI211_X1 _13299_ ( .A(_05797_ ), .B(_05736_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][17] ), .ZN(_05798_ ) );
AOI22_X1 _13300_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][17] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][17] ), .ZN(_05799_ ) );
AOI21_X1 _13301_ ( .A(_05747_ ), .B1(_05798_ ), .B2(_05799_ ), .ZN(_05800_ ) );
NOR2_X1 _13302_ ( .A1(_05796_ ), .A2(_05800_ ), .ZN(_05801_ ) );
NOR3_X1 _13303_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05801_ ), .ZN(_00388_ ) );
OR2_X1 _13304_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][16] ), .ZN(_05802_ ) );
OAI211_X1 _13305_ ( .A(_05802_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][16] ), .ZN(_05803_ ) );
AOI22_X1 _13306_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][16] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][16] ), .ZN(_05804_ ) );
AOI21_X1 _13307_ ( .A(fanout_net_8 ), .B1(_05803_ ), .B2(_05804_ ), .ZN(_05805_ ) );
OR2_X1 _13308_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][16] ), .ZN(_05806_ ) );
BUF_X4 _13309_ ( .A(_05724_ ), .Z(_05807_ ) );
OAI211_X1 _13310_ ( .A(_05806_ ), .B(_05807_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][16] ), .ZN(_05808_ ) );
AOI22_X1 _13311_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][16] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][16] ), .ZN(_05809_ ) );
AOI21_X1 _13312_ ( .A(_05747_ ), .B1(_05808_ ), .B2(_05809_ ), .ZN(_05810_ ) );
NOR2_X1 _13313_ ( .A1(_05805_ ), .A2(_05810_ ), .ZN(_05811_ ) );
NOR3_X1 _13314_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05811_ ), .ZN(_00389_ ) );
OR2_X1 _13315_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][15] ), .ZN(_05812_ ) );
OAI211_X1 _13316_ ( .A(_05812_ ), .B(_05725_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][15] ), .ZN(_05813_ ) );
AOI22_X1 _13317_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][15] ), .B1(_05731_ ), .B2(\u_icache.cblocks[3][15] ), .ZN(_05814_ ) );
AOI21_X1 _13318_ ( .A(fanout_net_8 ), .B1(_05813_ ), .B2(_05814_ ), .ZN(_05815_ ) );
OR2_X1 _13319_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][15] ), .ZN(_05816_ ) );
OAI211_X1 _13320_ ( .A(_05816_ ), .B(_05807_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][15] ), .ZN(_05817_ ) );
AOI22_X1 _13321_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][15] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][15] ), .ZN(_05818_ ) );
AOI21_X1 _13322_ ( .A(_05747_ ), .B1(_05817_ ), .B2(_05818_ ), .ZN(_05819_ ) );
NOR2_X1 _13323_ ( .A1(_05815_ ), .A2(_05819_ ), .ZN(_05820_ ) );
NOR3_X1 _13324_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05820_ ), .ZN(_00390_ ) );
OR2_X1 _13325_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][14] ), .ZN(_05821_ ) );
BUF_X4 _13326_ ( .A(_05724_ ), .Z(_05822_ ) );
OAI211_X1 _13327_ ( .A(_05821_ ), .B(_05822_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][14] ), .ZN(_05823_ ) );
BUF_X4 _13328_ ( .A(_05730_ ), .Z(_05824_ ) );
AOI22_X1 _13329_ ( .A1(_05728_ ), .A2(\u_icache.cblocks[2][14] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][14] ), .ZN(_05825_ ) );
AOI21_X1 _13330_ ( .A(fanout_net_8 ), .B1(_05823_ ), .B2(_05825_ ), .ZN(_05826_ ) );
OR2_X1 _13331_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][14] ), .ZN(_05827_ ) );
OAI211_X1 _13332_ ( .A(_05827_ ), .B(_05807_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][14] ), .ZN(_05828_ ) );
AOI22_X1 _13333_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][14] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][14] ), .ZN(_05829_ ) );
AOI21_X1 _13334_ ( .A(_05747_ ), .B1(_05828_ ), .B2(_05829_ ), .ZN(_05830_ ) );
NOR2_X1 _13335_ ( .A1(_05826_ ), .A2(_05830_ ), .ZN(_05831_ ) );
NOR3_X1 _13336_ ( .A1(_05718_ ), .A2(fanout_net_2 ), .A3(_05831_ ), .ZN(_00391_ ) );
BUF_X4 _13337_ ( .A(_00855_ ), .Z(_05832_ ) );
OR2_X1 _13338_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][13] ), .ZN(_05833_ ) );
OAI211_X1 _13339_ ( .A(_05833_ ), .B(_05822_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][13] ), .ZN(_05834_ ) );
BUF_X4 _13340_ ( .A(_05727_ ), .Z(_05835_ ) );
AOI22_X1 _13341_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][13] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][13] ), .ZN(_05836_ ) );
AOI21_X1 _13342_ ( .A(fanout_net_8 ), .B1(_05834_ ), .B2(_05836_ ), .ZN(_05837_ ) );
OR2_X1 _13343_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][13] ), .ZN(_05838_ ) );
OAI211_X1 _13344_ ( .A(_05838_ ), .B(_05807_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][13] ), .ZN(_05839_ ) );
AOI22_X1 _13345_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][13] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][13] ), .ZN(_05840_ ) );
AOI21_X1 _13346_ ( .A(_05747_ ), .B1(_05839_ ), .B2(_05840_ ), .ZN(_05841_ ) );
NOR2_X1 _13347_ ( .A1(_05837_ ), .A2(_05841_ ), .ZN(_05842_ ) );
NOR3_X1 _13348_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05842_ ), .ZN(_00392_ ) );
OR2_X1 _13349_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][12] ), .ZN(_05843_ ) );
OAI211_X1 _13350_ ( .A(_05843_ ), .B(_05822_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][12] ), .ZN(_05844_ ) );
AOI22_X1 _13351_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][12] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][12] ), .ZN(_05845_ ) );
AOI21_X1 _13352_ ( .A(fanout_net_8 ), .B1(_05844_ ), .B2(_05845_ ), .ZN(_05846_ ) );
BUF_X4 _13353_ ( .A(_05688_ ), .Z(_05847_ ) );
OR2_X1 _13354_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][12] ), .ZN(_05848_ ) );
OAI211_X1 _13355_ ( .A(_05848_ ), .B(_05807_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][12] ), .ZN(_05849_ ) );
AOI22_X1 _13356_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][12] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][12] ), .ZN(_05850_ ) );
AOI21_X1 _13357_ ( .A(_05847_ ), .B1(_05849_ ), .B2(_05850_ ), .ZN(_05851_ ) );
NOR2_X1 _13358_ ( .A1(_05846_ ), .A2(_05851_ ), .ZN(_05852_ ) );
NOR3_X1 _13359_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05852_ ), .ZN(_00393_ ) );
OR2_X1 _13360_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[5][29] ), .ZN(_05853_ ) );
OAI211_X1 _13361_ ( .A(_05853_ ), .B(_05822_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[4][29] ), .ZN(_05854_ ) );
AOI22_X1 _13362_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[6][29] ), .B1(_05824_ ), .B2(\u_icache.cblocks[7][29] ), .ZN(_05855_ ) );
AOI21_X1 _13363_ ( .A(_05690_ ), .B1(_05854_ ), .B2(_05855_ ), .ZN(_05856_ ) );
AOI22_X1 _13364_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[2][29] ), .B1(_05739_ ), .B2(\u_icache.cblocks[3][29] ), .ZN(_05857_ ) );
OR2_X1 _13365_ ( .A1(fanout_net_6 ), .A2(\u_icache.cblocks[0][29] ), .ZN(_05858_ ) );
OAI211_X1 _13366_ ( .A(_05858_ ), .B(_05724_ ), .C1(_05721_ ), .C2(\u_icache.cblocks[1][29] ), .ZN(_05859_ ) );
AOI21_X1 _13367_ ( .A(fanout_net_8 ), .B1(_05857_ ), .B2(_05859_ ), .ZN(_05860_ ) );
NOR2_X1 _13368_ ( .A1(_05856_ ), .A2(_05860_ ), .ZN(_05861_ ) );
NOR3_X1 _13369_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05861_ ), .ZN(_00394_ ) );
OR2_X1 _13370_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][11] ), .ZN(_05862_ ) );
OAI211_X1 _13371_ ( .A(_05862_ ), .B(_05822_ ), .C1(fanout_net_6 ), .C2(\u_icache.cblocks[0][11] ), .ZN(_05863_ ) );
AOI22_X1 _13372_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][11] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][11] ), .ZN(_05864_ ) );
AOI21_X1 _13373_ ( .A(fanout_net_8 ), .B1(_05863_ ), .B2(_05864_ ), .ZN(_05865_ ) );
OR2_X1 _13374_ ( .A1(_05766_ ), .A2(\u_icache.cblocks[5][11] ), .ZN(_05866_ ) );
OAI211_X1 _13375_ ( .A(_05866_ ), .B(_05807_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][11] ), .ZN(_05867_ ) );
AOI22_X1 _13376_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][11] ), .B1(_05769_ ), .B2(\u_icache.cblocks[7][11] ), .ZN(_05868_ ) );
AOI21_X1 _13377_ ( .A(_05847_ ), .B1(_05867_ ), .B2(_05868_ ), .ZN(_05869_ ) );
NOR2_X1 _13378_ ( .A1(_05865_ ), .A2(_05869_ ), .ZN(_05870_ ) );
NOR3_X1 _13379_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05870_ ), .ZN(_00395_ ) );
OR2_X1 _13380_ ( .A1(_05783_ ), .A2(\u_icache.cblocks[1][10] ), .ZN(_05871_ ) );
OAI211_X1 _13381_ ( .A(_05871_ ), .B(_05822_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][10] ), .ZN(_05872_ ) );
AOI22_X1 _13382_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][10] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][10] ), .ZN(_05873_ ) );
AOI21_X1 _13383_ ( .A(fanout_net_8 ), .B1(_05872_ ), .B2(_05873_ ), .ZN(_05874_ ) );
CLKBUF_X2 _13384_ ( .A(_05719_ ), .Z(_05875_ ) );
OR2_X1 _13385_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][10] ), .ZN(_05876_ ) );
OAI211_X1 _13386_ ( .A(_05876_ ), .B(_05807_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][10] ), .ZN(_05877_ ) );
BUF_X4 _13387_ ( .A(_05729_ ), .Z(_05878_ ) );
AOI22_X1 _13388_ ( .A1(_05779_ ), .A2(\u_icache.cblocks[6][10] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][10] ), .ZN(_05879_ ) );
AOI21_X1 _13389_ ( .A(_05847_ ), .B1(_05877_ ), .B2(_05879_ ), .ZN(_05880_ ) );
NOR2_X1 _13390_ ( .A1(_05874_ ), .A2(_05880_ ), .ZN(_05881_ ) );
NOR3_X1 _13391_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05881_ ), .ZN(_00396_ ) );
CLKBUF_X2 _13392_ ( .A(_05720_ ), .Z(_05882_ ) );
OR2_X1 _13393_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][9] ), .ZN(_05883_ ) );
OAI211_X1 _13394_ ( .A(_05883_ ), .B(_05822_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][9] ), .ZN(_05884_ ) );
AOI22_X1 _13395_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][9] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][9] ), .ZN(_05885_ ) );
AOI21_X1 _13396_ ( .A(fanout_net_8 ), .B1(_05884_ ), .B2(_05885_ ), .ZN(_05886_ ) );
OR2_X1 _13397_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][9] ), .ZN(_05887_ ) );
OAI211_X1 _13398_ ( .A(_05887_ ), .B(_05807_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][9] ), .ZN(_05888_ ) );
BUF_X4 _13399_ ( .A(_05727_ ), .Z(_05889_ ) );
AOI22_X1 _13400_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][9] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][9] ), .ZN(_05890_ ) );
AOI21_X1 _13401_ ( .A(_05847_ ), .B1(_05888_ ), .B2(_05890_ ), .ZN(_05891_ ) );
NOR2_X1 _13402_ ( .A1(_05886_ ), .A2(_05891_ ), .ZN(_05892_ ) );
NOR3_X1 _13403_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05892_ ), .ZN(_00397_ ) );
OR2_X1 _13404_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][8] ), .ZN(_05893_ ) );
OAI211_X1 _13405_ ( .A(_05893_ ), .B(_05822_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][8] ), .ZN(_05894_ ) );
AOI22_X1 _13406_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][8] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][8] ), .ZN(_05895_ ) );
AOI21_X1 _13407_ ( .A(fanout_net_8 ), .B1(_05894_ ), .B2(_05895_ ), .ZN(_05896_ ) );
OR2_X1 _13408_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][8] ), .ZN(_05897_ ) );
OAI211_X1 _13409_ ( .A(_05897_ ), .B(_05807_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][8] ), .ZN(_05898_ ) );
AOI22_X1 _13410_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][8] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][8] ), .ZN(_05899_ ) );
AOI21_X1 _13411_ ( .A(_05847_ ), .B1(_05898_ ), .B2(_05899_ ), .ZN(_05900_ ) );
NOR2_X1 _13412_ ( .A1(_05896_ ), .A2(_05900_ ), .ZN(_05901_ ) );
NOR3_X1 _13413_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05901_ ), .ZN(_00398_ ) );
OR2_X1 _13414_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][7] ), .ZN(_05902_ ) );
OAI211_X1 _13415_ ( .A(_05902_ ), .B(_05822_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][7] ), .ZN(_05903_ ) );
AOI22_X1 _13416_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][7] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][7] ), .ZN(_05904_ ) );
AOI21_X1 _13417_ ( .A(fanout_net_8 ), .B1(_05903_ ), .B2(_05904_ ), .ZN(_05905_ ) );
AOI22_X1 _13418_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[6][7] ), .B1(_05739_ ), .B2(\u_icache.cblocks[7][7] ), .ZN(_05906_ ) );
OR2_X1 _13419_ ( .A1(fanout_net_7 ), .A2(\u_icache.cblocks[4][7] ), .ZN(_05907_ ) );
OAI211_X1 _13420_ ( .A(_05907_ ), .B(_05724_ ), .C1(_05721_ ), .C2(\u_icache.cblocks[5][7] ), .ZN(_05908_ ) );
AOI21_X1 _13421_ ( .A(_05847_ ), .B1(_05906_ ), .B2(_05908_ ), .ZN(_05909_ ) );
NOR2_X1 _13422_ ( .A1(_05905_ ), .A2(_05909_ ), .ZN(_05910_ ) );
NOR3_X1 _13423_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05910_ ), .ZN(_00399_ ) );
OR2_X1 _13424_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][6] ), .ZN(_05911_ ) );
OAI211_X1 _13425_ ( .A(_05911_ ), .B(_05822_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][6] ), .ZN(_05912_ ) );
AOI22_X1 _13426_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][6] ), .B1(_05824_ ), .B2(\u_icache.cblocks[3][6] ), .ZN(_05913_ ) );
AOI21_X1 _13427_ ( .A(fanout_net_8 ), .B1(_05912_ ), .B2(_05913_ ), .ZN(_05914_ ) );
OR2_X1 _13428_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][6] ), .ZN(_05915_ ) );
OAI211_X1 _13429_ ( .A(_05915_ ), .B(_05807_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][6] ), .ZN(_05916_ ) );
AOI22_X1 _13430_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][6] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][6] ), .ZN(_05917_ ) );
AOI21_X1 _13431_ ( .A(_05847_ ), .B1(_05916_ ), .B2(_05917_ ), .ZN(_05918_ ) );
NOR2_X1 _13432_ ( .A1(_05914_ ), .A2(_05918_ ), .ZN(_05919_ ) );
NOR3_X1 _13433_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05919_ ), .ZN(_00400_ ) );
OR2_X1 _13434_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][5] ), .ZN(_05920_ ) );
BUF_X4 _13435_ ( .A(_05724_ ), .Z(_05921_ ) );
OAI211_X1 _13436_ ( .A(_05920_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][5] ), .ZN(_05922_ ) );
BUF_X4 _13437_ ( .A(_05730_ ), .Z(_05923_ ) );
AOI22_X1 _13438_ ( .A1(_05835_ ), .A2(\u_icache.cblocks[2][5] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][5] ), .ZN(_05924_ ) );
AOI21_X1 _13439_ ( .A(fanout_net_8 ), .B1(_05922_ ), .B2(_05924_ ), .ZN(_05925_ ) );
OR2_X1 _13440_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][5] ), .ZN(_05926_ ) );
BUF_X4 _13441_ ( .A(_05723_ ), .Z(_05927_ ) );
OAI211_X1 _13442_ ( .A(_05926_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][5] ), .ZN(_05928_ ) );
AOI22_X1 _13443_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][5] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][5] ), .ZN(_05929_ ) );
AOI21_X1 _13444_ ( .A(_05847_ ), .B1(_05928_ ), .B2(_05929_ ), .ZN(_05930_ ) );
NOR2_X1 _13445_ ( .A1(_05925_ ), .A2(_05930_ ), .ZN(_05931_ ) );
NOR3_X1 _13446_ ( .A1(_05832_ ), .A2(fanout_net_2 ), .A3(_05931_ ), .ZN(_00401_ ) );
BUF_X4 _13447_ ( .A(_00855_ ), .Z(_05932_ ) );
OR2_X1 _13448_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][4] ), .ZN(_05933_ ) );
OAI211_X1 _13449_ ( .A(_05933_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][4] ), .ZN(_05934_ ) );
BUF_X4 _13450_ ( .A(_05727_ ), .Z(_05935_ ) );
AOI22_X1 _13451_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][4] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][4] ), .ZN(_05936_ ) );
AOI21_X1 _13452_ ( .A(fanout_net_8 ), .B1(_05934_ ), .B2(_05936_ ), .ZN(_05937_ ) );
OR2_X1 _13453_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][4] ), .ZN(_05938_ ) );
OAI211_X1 _13454_ ( .A(_05938_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][4] ), .ZN(_05939_ ) );
AOI22_X1 _13455_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][4] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][4] ), .ZN(_05940_ ) );
AOI21_X1 _13456_ ( .A(_05847_ ), .B1(_05939_ ), .B2(_05940_ ), .ZN(_05941_ ) );
NOR2_X1 _13457_ ( .A1(_05937_ ), .A2(_05941_ ), .ZN(_05942_ ) );
NOR3_X1 _13458_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_05942_ ), .ZN(_00402_ ) );
OR2_X1 _13459_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][3] ), .ZN(_05943_ ) );
OAI211_X1 _13460_ ( .A(_05943_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][3] ), .ZN(_05944_ ) );
AOI22_X1 _13461_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][3] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][3] ), .ZN(_05945_ ) );
AOI21_X1 _13462_ ( .A(fanout_net_8 ), .B1(_05944_ ), .B2(_05945_ ), .ZN(_05946_ ) );
OR2_X1 _13463_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][3] ), .ZN(_05947_ ) );
OAI211_X1 _13464_ ( .A(_05947_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][3] ), .ZN(_05948_ ) );
AOI22_X1 _13465_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][3] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][3] ), .ZN(_05949_ ) );
AOI21_X1 _13466_ ( .A(_05847_ ), .B1(_05948_ ), .B2(_05949_ ), .ZN(_05950_ ) );
NOR2_X1 _13467_ ( .A1(_05946_ ), .A2(_05950_ ), .ZN(_05951_ ) );
NOR3_X1 _13468_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_05951_ ), .ZN(_00403_ ) );
OR2_X1 _13469_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][2] ), .ZN(_05952_ ) );
OAI211_X1 _13470_ ( .A(_05952_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][2] ), .ZN(_05953_ ) );
AOI22_X1 _13471_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][2] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][2] ), .ZN(_05954_ ) );
AOI21_X1 _13472_ ( .A(fanout_net_8 ), .B1(_05953_ ), .B2(_05954_ ), .ZN(_05955_ ) );
OR2_X1 _13473_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][2] ), .ZN(_05956_ ) );
OAI211_X1 _13474_ ( .A(_05956_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][2] ), .ZN(_05957_ ) );
AOI22_X1 _13475_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][2] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][2] ), .ZN(_05958_ ) );
AOI21_X1 _13476_ ( .A(_05689_ ), .B1(_05957_ ), .B2(_05958_ ), .ZN(_05959_ ) );
NOR2_X1 _13477_ ( .A1(_05955_ ), .A2(_05959_ ), .ZN(_05960_ ) );
NOR3_X1 _13478_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_05960_ ), .ZN(_00404_ ) );
OR2_X1 _13479_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][28] ), .ZN(_05961_ ) );
OAI211_X1 _13480_ ( .A(_05961_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][28] ), .ZN(_05962_ ) );
AOI22_X1 _13481_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][28] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][28] ), .ZN(_05963_ ) );
AOI21_X1 _13482_ ( .A(fanout_net_8 ), .B1(_05962_ ), .B2(_05963_ ), .ZN(_05964_ ) );
OR2_X1 _13483_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][28] ), .ZN(_05965_ ) );
OAI211_X1 _13484_ ( .A(_05965_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][28] ), .ZN(_05966_ ) );
AOI22_X1 _13485_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][28] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][28] ), .ZN(_05967_ ) );
AOI21_X1 _13486_ ( .A(_05689_ ), .B1(_05966_ ), .B2(_05967_ ), .ZN(_05968_ ) );
NOR2_X1 _13487_ ( .A1(_05964_ ), .A2(_05968_ ), .ZN(_05969_ ) );
NOR3_X1 _13488_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_05969_ ), .ZN(_00405_ ) );
OR2_X1 _13489_ ( .A1(_05882_ ), .A2(\u_icache.cblocks[1][1] ), .ZN(_05970_ ) );
OAI211_X1 _13490_ ( .A(_05970_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][1] ), .ZN(_05971_ ) );
AOI22_X1 _13491_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][1] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][1] ), .ZN(_05972_ ) );
AOI21_X1 _13492_ ( .A(fanout_net_8 ), .B1(_05971_ ), .B2(_05972_ ), .ZN(_05973_ ) );
OR2_X1 _13493_ ( .A1(_05875_ ), .A2(\u_icache.cblocks[5][1] ), .ZN(_05974_ ) );
OAI211_X1 _13494_ ( .A(_05974_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][1] ), .ZN(_05975_ ) );
AOI22_X1 _13495_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][1] ), .B1(_05878_ ), .B2(\u_icache.cblocks[7][1] ), .ZN(_05976_ ) );
AOI21_X1 _13496_ ( .A(_05689_ ), .B1(_05975_ ), .B2(_05976_ ), .ZN(_05977_ ) );
NOR2_X1 _13497_ ( .A1(_05973_ ), .A2(_05977_ ), .ZN(_05978_ ) );
NOR3_X1 _13498_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_05978_ ), .ZN(_00406_ ) );
OR2_X1 _13499_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[1][0] ), .ZN(_05979_ ) );
OAI211_X1 _13500_ ( .A(_05979_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][0] ), .ZN(_05980_ ) );
AOI22_X1 _13501_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][0] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][0] ), .ZN(_05981_ ) );
AOI21_X1 _13502_ ( .A(fanout_net_8 ), .B1(_05980_ ), .B2(_05981_ ), .ZN(_05982_ ) );
OR2_X1 _13503_ ( .A1(_05720_ ), .A2(\u_icache.cblocks[5][0] ), .ZN(_05983_ ) );
OAI211_X1 _13504_ ( .A(_05983_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][0] ), .ZN(_05984_ ) );
AOI22_X1 _13505_ ( .A1(_05889_ ), .A2(\u_icache.cblocks[6][0] ), .B1(_05730_ ), .B2(\u_icache.cblocks[7][0] ), .ZN(_05985_ ) );
AOI21_X1 _13506_ ( .A(_05689_ ), .B1(_05984_ ), .B2(_05985_ ), .ZN(_05986_ ) );
NOR2_X1 _13507_ ( .A1(_05982_ ), .A2(_05986_ ), .ZN(_05987_ ) );
NOR3_X1 _13508_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_05987_ ), .ZN(_00407_ ) );
OR2_X1 _13509_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[1][27] ), .ZN(_05988_ ) );
OAI211_X1 _13510_ ( .A(_05988_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][27] ), .ZN(_05989_ ) );
AOI22_X1 _13511_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][27] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][27] ), .ZN(_05990_ ) );
AOI21_X1 _13512_ ( .A(fanout_net_8 ), .B1(_05989_ ), .B2(_05990_ ), .ZN(_05991_ ) );
OR2_X1 _13513_ ( .A1(_05720_ ), .A2(\u_icache.cblocks[5][27] ), .ZN(_05992_ ) );
OAI211_X1 _13514_ ( .A(_05992_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][27] ), .ZN(_05993_ ) );
AOI22_X1 _13515_ ( .A1(_05727_ ), .A2(\u_icache.cblocks[6][27] ), .B1(_05730_ ), .B2(\u_icache.cblocks[7][27] ), .ZN(_05994_ ) );
AOI21_X1 _13516_ ( .A(_05689_ ), .B1(_05993_ ), .B2(_05994_ ), .ZN(_05995_ ) );
NOR2_X1 _13517_ ( .A1(_05991_ ), .A2(_05995_ ), .ZN(_05996_ ) );
NOR3_X1 _13518_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_05996_ ), .ZN(_00408_ ) );
OR2_X1 _13519_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[1][26] ), .ZN(_05997_ ) );
OAI211_X1 _13520_ ( .A(_05997_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[0][26] ), .ZN(_05998_ ) );
AOI22_X1 _13521_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][26] ), .B1(_05923_ ), .B2(\u_icache.cblocks[3][26] ), .ZN(_05999_ ) );
AOI21_X1 _13522_ ( .A(fanout_net_8 ), .B1(_05998_ ), .B2(_05999_ ), .ZN(_06000_ ) );
OR2_X1 _13523_ ( .A1(_05720_ ), .A2(\u_icache.cblocks[5][26] ), .ZN(_06001_ ) );
OAI211_X1 _13524_ ( .A(_06001_ ), .B(_05927_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][26] ), .ZN(_06002_ ) );
AOI22_X1 _13525_ ( .A1(_05727_ ), .A2(\u_icache.cblocks[6][26] ), .B1(_05730_ ), .B2(\u_icache.cblocks[7][26] ), .ZN(_06003_ ) );
AOI21_X1 _13526_ ( .A(_05689_ ), .B1(_06002_ ), .B2(_06003_ ), .ZN(_06004_ ) );
NOR2_X1 _13527_ ( .A1(_06000_ ), .A2(_06004_ ), .ZN(_06005_ ) );
NOR3_X1 _13528_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_06005_ ), .ZN(_00409_ ) );
OR2_X1 _13529_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[5][25] ), .ZN(_06006_ ) );
OAI211_X1 _13530_ ( .A(_06006_ ), .B(_05921_ ), .C1(fanout_net_7 ), .C2(\u_icache.cblocks[4][25] ), .ZN(_06007_ ) );
AOI22_X1 _13531_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[6][25] ), .B1(_05923_ ), .B2(\u_icache.cblocks[7][25] ), .ZN(_06008_ ) );
AOI21_X1 _13532_ ( .A(_05690_ ), .B1(_06007_ ), .B2(_06008_ ), .ZN(_06009_ ) );
AOI22_X1 _13533_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[2][25] ), .B1(_05739_ ), .B2(\u_icache.cblocks[3][25] ), .ZN(_06010_ ) );
OR2_X1 _13534_ ( .A1(\fc_addr [2] ), .A2(\u_icache.cblocks[0][25] ), .ZN(_06011_ ) );
OAI211_X1 _13535_ ( .A(_06011_ ), .B(_05724_ ), .C1(_05721_ ), .C2(\u_icache.cblocks[1][25] ), .ZN(_06012_ ) );
AOI21_X1 _13536_ ( .A(\fc_addr [4] ), .B1(_06010_ ), .B2(_06012_ ), .ZN(_06013_ ) );
NOR2_X1 _13537_ ( .A1(_06009_ ), .A2(_06013_ ), .ZN(_06014_ ) );
NOR3_X1 _13538_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_06014_ ), .ZN(_00410_ ) );
OR2_X1 _13539_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[1][24] ), .ZN(_06015_ ) );
OAI211_X1 _13540_ ( .A(_06015_ ), .B(_05736_ ), .C1(\fc_addr [2] ), .C2(\u_icache.cblocks[0][24] ), .ZN(_06016_ ) );
AOI22_X1 _13541_ ( .A1(_05935_ ), .A2(\u_icache.cblocks[2][24] ), .B1(_05739_ ), .B2(\u_icache.cblocks[3][24] ), .ZN(_06017_ ) );
AOI21_X1 _13542_ ( .A(\fc_addr [4] ), .B1(_06016_ ), .B2(_06017_ ), .ZN(_06018_ ) );
OR2_X1 _13543_ ( .A1(_05720_ ), .A2(\u_icache.cblocks[5][24] ), .ZN(_06019_ ) );
OAI211_X1 _13544_ ( .A(_06019_ ), .B(_05927_ ), .C1(\fc_addr [2] ), .C2(\u_icache.cblocks[4][24] ), .ZN(_06020_ ) );
AOI22_X1 _13545_ ( .A1(_05727_ ), .A2(\u_icache.cblocks[6][24] ), .B1(_05730_ ), .B2(\u_icache.cblocks[7][24] ), .ZN(_06021_ ) );
AOI21_X1 _13546_ ( .A(_05689_ ), .B1(_06020_ ), .B2(_06021_ ), .ZN(_06022_ ) );
NOR2_X1 _13547_ ( .A1(_06018_ ), .A2(_06022_ ), .ZN(_06023_ ) );
NOR3_X1 _13548_ ( .A1(_05932_ ), .A2(fanout_net_3 ), .A3(_06023_ ), .ZN(_00411_ ) );
OR2_X1 _13549_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[5][23] ), .ZN(_06024_ ) );
OAI211_X1 _13550_ ( .A(_06024_ ), .B(_05736_ ), .C1(\fc_addr [2] ), .C2(\u_icache.cblocks[4][23] ), .ZN(_06025_ ) );
AOI22_X1 _13551_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[6][23] ), .B1(_05739_ ), .B2(\u_icache.cblocks[7][23] ), .ZN(_06026_ ) );
AOI21_X1 _13552_ ( .A(_05690_ ), .B1(_06025_ ), .B2(_06026_ ), .ZN(_06027_ ) );
AOI22_X1 _13553_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[2][23] ), .B1(_05739_ ), .B2(\u_icache.cblocks[3][23] ), .ZN(_06028_ ) );
OR2_X1 _13554_ ( .A1(\fc_addr [2] ), .A2(\u_icache.cblocks[0][23] ), .ZN(_06029_ ) );
OAI211_X1 _13555_ ( .A(_06029_ ), .B(_05724_ ), .C1(_05721_ ), .C2(\u_icache.cblocks[1][23] ), .ZN(_06030_ ) );
AOI21_X1 _13556_ ( .A(\fc_addr [4] ), .B1(_06028_ ), .B2(_06030_ ), .ZN(_06031_ ) );
NOR2_X1 _13557_ ( .A1(_06027_ ), .A2(_06031_ ), .ZN(_06032_ ) );
NOR3_X1 _13558_ ( .A1(_00856_ ), .A2(fanout_net_3 ), .A3(_06032_ ), .ZN(_00412_ ) );
OR2_X1 _13559_ ( .A1(_05734_ ), .A2(\u_icache.cblocks[1][22] ), .ZN(_06033_ ) );
OAI211_X1 _13560_ ( .A(_06033_ ), .B(_05736_ ), .C1(\fc_addr [2] ), .C2(\u_icache.cblocks[0][22] ), .ZN(_06034_ ) );
AOI22_X1 _13561_ ( .A1(_05738_ ), .A2(\u_icache.cblocks[2][22] ), .B1(_05739_ ), .B2(\u_icache.cblocks[3][22] ), .ZN(_06035_ ) );
AOI21_X1 _13562_ ( .A(\fc_addr [4] ), .B1(_06034_ ), .B2(_06035_ ), .ZN(_06036_ ) );
OR2_X1 _13563_ ( .A1(_05720_ ), .A2(\u_icache.cblocks[5][22] ), .ZN(_06037_ ) );
OAI211_X1 _13564_ ( .A(_06037_ ), .B(_05724_ ), .C1(\fc_addr [2] ), .C2(\u_icache.cblocks[4][22] ), .ZN(_06038_ ) );
AOI22_X1 _13565_ ( .A1(_05727_ ), .A2(\u_icache.cblocks[6][22] ), .B1(_05730_ ), .B2(\u_icache.cblocks[7][22] ), .ZN(_06039_ ) );
AOI21_X1 _13566_ ( .A(_05689_ ), .B1(_06038_ ), .B2(_06039_ ), .ZN(_06040_ ) );
NOR2_X1 _13567_ ( .A1(_06036_ ), .A2(_06040_ ), .ZN(_06041_ ) );
NOR3_X1 _13568_ ( .A1(_00856_ ), .A2(fanout_net_3 ), .A3(_06041_ ), .ZN(_00413_ ) );
AND2_X1 _13569_ ( .A1(\u_icache.count [1] ), .A2(\u_icache.count [0] ), .ZN(_06042_ ) );
INV_X1 _13570_ ( .A(\u_icache.count [2] ), .ZN(_06043_ ) );
XNOR2_X1 _13571_ ( .A(_06042_ ), .B(_06043_ ), .ZN(_06044_ ) );
AND4_X1 _13572_ ( .A1(_00863_ ), .A2(_05550_ ), .A3(_05551_ ), .A4(_06044_ ), .ZN(_00415_ ) );
INV_X1 _13573_ ( .A(_05640_ ), .ZN(_06045_ ) );
NOR2_X1 _13574_ ( .A1(\u_icache.count [1] ), .A2(\u_icache.count [0] ), .ZN(_06046_ ) );
NOR4_X1 _13575_ ( .A1(_06045_ ), .A2(_05548_ ), .A3(_06042_ ), .A4(_06046_ ), .ZN(_00416_ ) );
INV_X1 _13576_ ( .A(_05550_ ), .ZN(_06047_ ) );
BUF_X4 _13577_ ( .A(_01149_ ), .Z(_06048_ ) );
NOR4_X1 _13578_ ( .A1(_06047_ ), .A2(\u_icache.count [0] ), .A3(_05548_ ), .A4(_06048_ ), .ZN(_00417_ ) );
INV_X1 _13579_ ( .A(ifu_ready ), .ZN(_06049_ ) );
AND3_X1 _13580_ ( .A1(_05481_ ), .A2(_05545_ ), .A3(_06049_ ), .ZN(_06050_ ) );
OAI21_X1 _13581_ ( .A(_06050_ ), .B1(_05400_ ), .B2(_05402_ ), .ZN(_06051_ ) );
AND2_X1 _13582_ ( .A1(_06046_ ), .A2(\u_icache.count [2] ), .ZN(\u_icache.cvalids_$_SDFFE_PP0P__Q_E ) );
INV_X1 _13583_ ( .A(\u_icache.cvalids_$_SDFFE_PP0P__Q_E ), .ZN(_06052_ ) );
NAND2_X1 _13584_ ( .A1(_06051_ ), .A2(_06052_ ), .ZN(\u_icache.cready_$_ANDNOT__B_Y_$_OR__B_Y ) );
AOI21_X1 _13585_ ( .A(_04462_ ), .B1(_06051_ ), .B2(_06052_ ), .ZN(_00418_ ) );
AOI211_X1 _13586_ ( .A(fanout_net_3 ), .B(_00882_ ), .C1(_05690_ ), .C2(_05484_ ), .ZN(_00419_ ) );
AOI211_X1 _13587_ ( .A(fanout_net_3 ), .B(_00882_ ), .C1(\fc_addr [4] ), .C2(_05483_ ), .ZN(_00420_ ) );
AND4_X1 _13588_ ( .A1(_06043_ ), .A2(icah_ready ), .A3(_04476_ ), .A4(_06042_ ), .ZN(_00421_ ) );
BUF_X2 _13589_ ( .A(_00770_ ), .Z(\u_ifu.inst_ok_$_ANDNOT__A_Y ) );
INV_X2 _13590_ ( .A(_00769_ ), .ZN(_06053_ ) );
BUF_X4 _13591_ ( .A(_06053_ ), .Z(_06054_ ) );
BUF_X4 _13592_ ( .A(_06054_ ), .Z(_06055_ ) );
NOR4_X1 _13593_ ( .A1(_04466_ ), .A2(fanout_net_3 ), .A3(_04467_ ), .A4(_06055_ ), .ZN(_00422_ ) );
AND3_X1 _13594_ ( .A1(_04465_ ), .A2(\fd_inst [31] ), .A3(_04468_ ), .ZN(_00423_ ) );
AND3_X1 _13595_ ( .A1(_04465_ ), .A2(\fd_inst [30] ), .A3(_04468_ ), .ZN(_00424_ ) );
CLKBUF_X2 _13596_ ( .A(_00862_ ), .Z(_06056_ ) );
AND3_X1 _13597_ ( .A1(_06056_ ), .A2(\fd_inst [21] ), .A3(_04468_ ), .ZN(_00425_ ) );
AND3_X1 _13598_ ( .A1(_06056_ ), .A2(\fd_inst [20] ), .A3(_04468_ ), .ZN(_00426_ ) );
AND3_X1 _13599_ ( .A1(_06056_ ), .A2(\fd_inst [19] ), .A3(_04468_ ), .ZN(_00427_ ) );
AND3_X1 _13600_ ( .A1(_06056_ ), .A2(\fd_inst [18] ), .A3(_04468_ ), .ZN(_00428_ ) );
AND3_X1 _13601_ ( .A1(_06056_ ), .A2(\fd_inst [17] ), .A3(_04468_ ), .ZN(_00429_ ) );
AND3_X1 _13602_ ( .A1(_06056_ ), .A2(\fd_inst [16] ), .A3(_04468_ ), .ZN(_00430_ ) );
AND3_X1 _13603_ ( .A1(_06056_ ), .A2(\fd_inst [15] ), .A3(_04468_ ), .ZN(_00431_ ) );
CLKBUF_X2 _13604_ ( .A(_00865_ ), .Z(_06057_ ) );
AND3_X1 _13605_ ( .A1(_06056_ ), .A2(\fd_inst [14] ), .A3(_06057_ ), .ZN(_00432_ ) );
AND3_X1 _13606_ ( .A1(_06056_ ), .A2(\fd_inst [13] ), .A3(_06057_ ), .ZN(_00433_ ) );
AND3_X1 _13607_ ( .A1(_06056_ ), .A2(\fd_inst [12] ), .A3(_06057_ ), .ZN(_00434_ ) );
CLKBUF_X2 _13608_ ( .A(_00862_ ), .Z(_06058_ ) );
AND3_X1 _13609_ ( .A1(_06058_ ), .A2(\fd_inst [29] ), .A3(_06057_ ), .ZN(_00435_ ) );
AND3_X1 _13610_ ( .A1(_06058_ ), .A2(\fd_inst [11] ), .A3(_06057_ ), .ZN(_00436_ ) );
AND3_X1 _13611_ ( .A1(_06058_ ), .A2(\fd_inst [10] ), .A3(_06057_ ), .ZN(_00437_ ) );
AND3_X1 _13612_ ( .A1(_06058_ ), .A2(\fd_inst [9] ), .A3(_06057_ ), .ZN(_00438_ ) );
AND3_X1 _13613_ ( .A1(_06058_ ), .A2(\fd_inst [8] ), .A3(_06057_ ), .ZN(_00439_ ) );
AND3_X1 _13614_ ( .A1(_06058_ ), .A2(\fd_inst [7] ), .A3(_06057_ ), .ZN(_00440_ ) );
AND3_X1 _13615_ ( .A1(_06058_ ), .A2(\fd_inst [6] ), .A3(_06057_ ), .ZN(_00441_ ) );
CLKBUF_X2 _13616_ ( .A(_00865_ ), .Z(_06059_ ) );
AND3_X1 _13617_ ( .A1(_06058_ ), .A2(\fd_inst [5] ), .A3(_06059_ ), .ZN(_00442_ ) );
AND3_X1 _13618_ ( .A1(_06058_ ), .A2(\fd_inst [4] ), .A3(_06059_ ), .ZN(_00443_ ) );
AND3_X1 _13619_ ( .A1(_06058_ ), .A2(\fd_inst [3] ), .A3(_06059_ ), .ZN(_00444_ ) );
CLKBUF_X2 _13620_ ( .A(_00862_ ), .Z(_06060_ ) );
AND3_X1 _13621_ ( .A1(_06060_ ), .A2(\fd_inst [2] ), .A3(_06059_ ), .ZN(_00445_ ) );
AND3_X1 _13622_ ( .A1(_06060_ ), .A2(\fd_inst [28] ), .A3(_06059_ ), .ZN(_00446_ ) );
AND3_X1 _13623_ ( .A1(_06060_ ), .A2(\fd_inst [1] ), .A3(_06059_ ), .ZN(_00447_ ) );
AND3_X1 _13624_ ( .A1(_06060_ ), .A2(\fd_inst [0] ), .A3(_06059_ ), .ZN(_00448_ ) );
AND3_X1 _13625_ ( .A1(_06060_ ), .A2(\fd_inst [27] ), .A3(_06059_ ), .ZN(_00449_ ) );
AND3_X1 _13626_ ( .A1(_06060_ ), .A2(\fd_inst [26] ), .A3(_06059_ ), .ZN(_00450_ ) );
AND3_X1 _13627_ ( .A1(_06060_ ), .A2(\fd_inst [25] ), .A3(_06059_ ), .ZN(_00451_ ) );
CLKBUF_X2 _13628_ ( .A(_00865_ ), .Z(_06061_ ) );
AND3_X1 _13629_ ( .A1(_06060_ ), .A2(\fd_inst [24] ), .A3(_06061_ ), .ZN(_00452_ ) );
AND3_X1 _13630_ ( .A1(_06060_ ), .A2(\fd_inst [23] ), .A3(_06061_ ), .ZN(_00453_ ) );
AND3_X1 _13631_ ( .A1(_06060_ ), .A2(\fd_inst [22] ), .A3(_06061_ ), .ZN(_00454_ ) );
NOR4_X1 _13632_ ( .A1(_04466_ ), .A2(fanout_net_3 ), .A3(_04467_ ), .A4(_05442_ ), .ZN(_00455_ ) );
BUF_X4 _13633_ ( .A(_00855_ ), .Z(_06062_ ) );
NOR4_X1 _13634_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_04467_ ), .A4(_05525_ ), .ZN(_00456_ ) );
NOR4_X1 _13635_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_04467_ ), .A4(_05650_ ), .ZN(_00457_ ) );
NOR4_X1 _13636_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_04467_ ), .A4(_05530_ ), .ZN(_00458_ ) );
NOR4_X1 _13637_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_04467_ ), .A4(_05654_ ), .ZN(_00459_ ) );
NOR4_X1 _13638_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_04467_ ), .A4(_05540_ ), .ZN(_00460_ ) );
BUF_X4 _13639_ ( .A(_00858_ ), .Z(_06063_ ) );
NOR4_X1 _13640_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05657_ ), .ZN(_00461_ ) );
NOR4_X1 _13641_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05439_ ), .ZN(_00462_ ) );
NOR4_X1 _13642_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05661_ ), .ZN(_00463_ ) );
NOR4_X1 _13643_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05664_ ), .ZN(_00464_ ) );
NOR4_X1 _13644_ ( .A1(_06062_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05425_ ), .ZN(_00465_ ) );
BUF_X4 _13645_ ( .A(_00855_ ), .Z(_06064_ ) );
NOR4_X1 _13646_ ( .A1(_06064_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05516_ ), .ZN(_00466_ ) );
NOR4_X1 _13647_ ( .A1(_06064_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05416_ ), .ZN(_00467_ ) );
NOR4_X1 _13648_ ( .A1(_06064_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05533_ ), .ZN(_00468_ ) );
NOR4_X1 _13649_ ( .A1(_06064_ ), .A2(fanout_net_3 ), .A3(_06063_ ), .A4(_05676_ ), .ZN(_00469_ ) );
NOR4_X1 _13650_ ( .A1(_06064_ ), .A2(fanout_net_4 ), .A3(_06063_ ), .A4(_05678_ ), .ZN(_00470_ ) );
BUF_X4 _13651_ ( .A(_00858_ ), .Z(_06065_ ) );
NOR4_X1 _13652_ ( .A1(_06064_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05497_ ), .ZN(_00471_ ) );
NOR4_X1 _13653_ ( .A1(_06064_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05681_ ), .ZN(_00472_ ) );
NOR4_X1 _13654_ ( .A1(_06064_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05487_ ), .ZN(_00473_ ) );
NOR4_X1 _13655_ ( .A1(_06064_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05685_ ), .ZN(_00474_ ) );
NOR4_X1 _13656_ ( .A1(_06064_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05690_ ), .ZN(_00475_ ) );
BUF_X4 _13657_ ( .A(_00855_ ), .Z(_06066_ ) );
NOR4_X1 _13658_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05725_ ), .ZN(_00476_ ) );
NOR4_X1 _13659_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05721_ ), .ZN(_00477_ ) );
NOR4_X1 _13660_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05693_ ), .ZN(_00478_ ) );
AND3_X1 _13661_ ( .A1(_04454_ ), .A2(\fc_addr [1] ), .A3(_06061_ ), .ZN(_00479_ ) );
AND3_X1 _13662_ ( .A1(_04454_ ), .A2(\fc_addr [0] ), .A3(_06061_ ), .ZN(_00480_ ) );
NOR4_X1 _13663_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05462_ ), .ZN(_00481_ ) );
NOR4_X1 _13664_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06065_ ), .A4(_05469_ ), .ZN(_00482_ ) );
BUF_X4 _13665_ ( .A(_00858_ ), .Z(_06067_ ) );
NOR4_X1 _13666_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06067_ ), .A4(_05458_ ), .ZN(_00483_ ) );
NOR4_X1 _13667_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06067_ ), .A4(_05708_ ), .ZN(_00484_ ) );
NOR4_X1 _13668_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06067_ ), .A4(_05476_ ), .ZN(_00485_ ) );
NOR4_X1 _13669_ ( .A1(_06066_ ), .A2(fanout_net_4 ), .A3(_06067_ ), .A4(_05451_ ), .ZN(_00486_ ) );
BUF_X2 _13670_ ( .A(_00640_ ), .Z(_06068_ ) );
BUF_X2 _13671_ ( .A(_06068_ ), .Z(_06069_ ) );
AND3_X1 _13672_ ( .A1(_06069_ ), .A2(_00829_ ), .A3(\cf_inst [31] ), .ZN(_00487_ ) );
CLKBUF_X2 _13673_ ( .A(_06068_ ), .Z(_06070_ ) );
AND3_X1 _13674_ ( .A1(_06070_ ), .A2(_00829_ ), .A3(\cf_inst [30] ), .ZN(_00488_ ) );
AND3_X1 _13675_ ( .A1(_06070_ ), .A2(_00829_ ), .A3(\cf_inst [21] ), .ZN(_00489_ ) );
AND3_X1 _13676_ ( .A1(_06070_ ), .A2(_00829_ ), .A3(\cf_inst [20] ), .ZN(_00490_ ) );
CLKBUF_X2 _13677_ ( .A(_00771_ ), .Z(_06071_ ) );
AND3_X1 _13678_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(\cf_inst [19] ), .ZN(_00491_ ) );
AND3_X1 _13679_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(\cf_inst [18] ), .ZN(_00492_ ) );
AND3_X1 _13680_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(\cf_inst [17] ), .ZN(_00493_ ) );
AND3_X1 _13681_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(\cf_inst [16] ), .ZN(_00494_ ) );
AND3_X1 _13682_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(\cf_inst [15] ), .ZN(_00495_ ) );
AND3_X1 _13683_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(\cf_inst [14] ), .ZN(_00496_ ) );
AND3_X1 _13684_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(\cf_inst [13] ), .ZN(_00497_ ) );
CLKBUF_X2 _13685_ ( .A(_00865_ ), .Z(_06072_ ) );
AND3_X1 _13686_ ( .A1(_06072_ ), .A2(_06071_ ), .A3(\cf_inst [12] ), .ZN(_00498_ ) );
AND3_X1 _13687_ ( .A1(_06072_ ), .A2(_06071_ ), .A3(\cf_inst [29] ), .ZN(_00499_ ) );
AND3_X1 _13688_ ( .A1(_06072_ ), .A2(_06071_ ), .A3(\cf_inst [11] ), .ZN(_00500_ ) );
CLKBUF_X2 _13689_ ( .A(_00771_ ), .Z(_06073_ ) );
AND3_X1 _13690_ ( .A1(_06072_ ), .A2(_06073_ ), .A3(\cf_inst [10] ), .ZN(_00501_ ) );
AND3_X1 _13691_ ( .A1(_06072_ ), .A2(_06073_ ), .A3(\cf_inst [9] ), .ZN(_00502_ ) );
AND3_X1 _13692_ ( .A1(_06072_ ), .A2(_06073_ ), .A3(\cf_inst [8] ), .ZN(_00503_ ) );
AND3_X1 _13693_ ( .A1(_06072_ ), .A2(_06073_ ), .A3(\cf_inst [7] ), .ZN(_00504_ ) );
AND3_X1 _13694_ ( .A1(_06072_ ), .A2(_06073_ ), .A3(\cf_inst [6] ), .ZN(_00505_ ) );
AND3_X1 _13695_ ( .A1(_06072_ ), .A2(_06073_ ), .A3(\cf_inst [5] ), .ZN(_00506_ ) );
AND3_X1 _13696_ ( .A1(_06072_ ), .A2(_06073_ ), .A3(\cf_inst [4] ), .ZN(_00507_ ) );
CLKBUF_X2 _13697_ ( .A(_00865_ ), .Z(_06074_ ) );
AND3_X1 _13698_ ( .A1(_06074_ ), .A2(_06073_ ), .A3(\cf_inst [3] ), .ZN(_00508_ ) );
AND3_X1 _13699_ ( .A1(_06074_ ), .A2(_06073_ ), .A3(\cf_inst [2] ), .ZN(_00509_ ) );
AND3_X1 _13700_ ( .A1(_06074_ ), .A2(_06073_ ), .A3(\cf_inst [28] ), .ZN(_00510_ ) );
AND3_X1 _13701_ ( .A1(_06074_ ), .A2(_00778_ ), .A3(\cf_inst [1] ), .ZN(_00511_ ) );
AND3_X1 _13702_ ( .A1(_06074_ ), .A2(_00778_ ), .A3(\cf_inst [0] ), .ZN(_00512_ ) );
AND3_X1 _13703_ ( .A1(_06074_ ), .A2(_00778_ ), .A3(\cf_inst [27] ), .ZN(_00513_ ) );
AND3_X1 _13704_ ( .A1(_06074_ ), .A2(_00778_ ), .A3(\cf_inst [26] ), .ZN(_00514_ ) );
AND3_X1 _13705_ ( .A1(_06074_ ), .A2(_00778_ ), .A3(\cf_inst [25] ), .ZN(_00515_ ) );
AND3_X1 _13706_ ( .A1(_06074_ ), .A2(_00778_ ), .A3(\cf_inst [24] ), .ZN(_00516_ ) );
AND3_X1 _13707_ ( .A1(_06074_ ), .A2(_00778_ ), .A3(\cf_inst [23] ), .ZN(_00517_ ) );
AND3_X1 _13708_ ( .A1(_00866_ ), .A2(_00778_ ), .A3(\cf_inst [22] ), .ZN(_00518_ ) );
NOR2_X1 _13709_ ( .A1(_05403_ ), .A2(_06049_ ), .ZN(\u_icache.cready_$_ANDNOT__A_Y ) );
NOR3_X1 _13710_ ( .A1(_05403_ ), .A2(_06049_ ), .A3(_04455_ ), .ZN(_00519_ ) );
AOI211_X1 _13711_ ( .A(_00765_ ), .B(_00880_ ), .C1(_00746_ ), .C2(_00758_ ), .ZN(_00520_ ) );
AND3_X1 _13712_ ( .A1(_01595_ ), .A2(_00858_ ), .A3(_01598_ ), .ZN(_06075_ ) );
NAND3_X4 _13713_ ( .A1(\fc_addr [5] ), .A2(\fc_addr [3] ), .A3(\fc_addr [2] ), .ZN(_06076_ ) );
NOR2_X1 _13714_ ( .A1(_06076_ ), .A2(_05688_ ), .ZN(_06077_ ) );
AND2_X2 _13715_ ( .A1(_06077_ ), .A2(\fc_addr [6] ), .ZN(_06078_ ) );
AND2_X2 _13716_ ( .A1(_06078_ ), .A2(\fc_addr [7] ), .ZN(_06079_ ) );
AND2_X2 _13717_ ( .A1(_06079_ ), .A2(\fc_addr [8] ), .ZN(_06080_ ) );
AND2_X4 _13718_ ( .A1(_06080_ ), .A2(\fc_addr [9] ), .ZN(_06081_ ) );
AND2_X4 _13719_ ( .A1(_06081_ ), .A2(\fc_addr [10] ), .ZN(_06082_ ) );
AND3_X4 _13720_ ( .A1(_06082_ ), .A2(\fc_addr [12] ), .A3(\fc_addr [11] ), .ZN(_06083_ ) );
AND2_X1 _13721_ ( .A1(_06083_ ), .A2(\fc_addr [13] ), .ZN(_06084_ ) );
AND2_X2 _13722_ ( .A1(_06084_ ), .A2(\fc_addr [14] ), .ZN(_06085_ ) );
AND2_X4 _13723_ ( .A1(_06085_ ), .A2(\fc_addr [15] ), .ZN(_06086_ ) );
AND2_X2 _13724_ ( .A1(_06086_ ), .A2(\fc_addr [16] ), .ZN(_06087_ ) );
AND2_X2 _13725_ ( .A1(_06087_ ), .A2(\fc_addr [17] ), .ZN(_06088_ ) );
AND2_X1 _13726_ ( .A1(_06088_ ), .A2(\fc_addr [18] ), .ZN(_06089_ ) );
AND2_X1 _13727_ ( .A1(_06089_ ), .A2(\fc_addr [19] ), .ZN(_06090_ ) );
AND3_X2 _13728_ ( .A1(_06090_ ), .A2(\fc_addr [21] ), .A3(\fc_addr [20] ), .ZN(_06091_ ) );
AND3_X1 _13729_ ( .A1(_06091_ ), .A2(\fc_addr [23] ), .A3(\fc_addr [22] ), .ZN(_06092_ ) );
AND3_X2 _13730_ ( .A1(_06092_ ), .A2(\fc_addr [25] ), .A3(\fc_addr [24] ), .ZN(_06093_ ) );
AND3_X2 _13731_ ( .A1(_06093_ ), .A2(\fc_addr [27] ), .A3(\fc_addr [26] ), .ZN(_06094_ ) );
NAND3_X2 _13732_ ( .A1(_06094_ ), .A2(\fc_addr [29] ), .A3(\fc_addr [28] ), .ZN(_06095_ ) );
XNOR2_X1 _13733_ ( .A(_06095_ ), .B(_05525_ ), .ZN(_06096_ ) );
MUX2_X2 _13734_ ( .A(_06096_ ), .B(_04654_ ), .S(_06054_ ), .Z(_06097_ ) );
AOI211_X1 _13735_ ( .A(fanout_net_4 ), .B(_06075_ ), .C1(_06097_ ), .C2(_06069_ ), .ZN(_00521_ ) );
AND3_X1 _13736_ ( .A1(_02171_ ), .A2(_00858_ ), .A3(_02172_ ), .ZN(_06098_ ) );
NAND4_X1 _13737_ ( .A1(\fc_addr [17] ), .A2(\fc_addr [16] ), .A3(\fc_addr [15] ), .A4(\fc_addr [14] ), .ZN(_06099_ ) );
NAND2_X1 _13738_ ( .A1(\fc_addr [11] ), .A2(\fc_addr [10] ), .ZN(_06100_ ) );
NOR4_X1 _13739_ ( .A1(_06099_ ), .A2(_06100_ ), .A3(_05425_ ), .A4(_05516_ ), .ZN(_06101_ ) );
AND2_X2 _13740_ ( .A1(_06081_ ), .A2(_06101_ ), .ZN(_06102_ ) );
AND4_X1 _13741_ ( .A1(\fc_addr [25] ), .A2(\fc_addr [24] ), .A3(\fc_addr [23] ), .A4(\fc_addr [22] ), .ZN(_06103_ ) );
AND2_X1 _13742_ ( .A1(\fc_addr [19] ), .A2(\fc_addr [18] ), .ZN(_06104_ ) );
AND4_X1 _13743_ ( .A1(\fc_addr [21] ), .A2(_06103_ ), .A3(\fc_addr [20] ), .A4(_06104_ ), .ZN(_06105_ ) );
AND2_X1 _13744_ ( .A1(_06102_ ), .A2(_06105_ ), .ZN(_06106_ ) );
AND3_X1 _13745_ ( .A1(_06106_ ), .A2(\fc_addr [27] ), .A3(\fc_addr [26] ), .ZN(_06107_ ) );
NAND2_X1 _13746_ ( .A1(_06107_ ), .A2(\fc_addr [28] ), .ZN(_06108_ ) );
NAND2_X1 _13747_ ( .A1(_06108_ ), .A2(\fc_addr [29] ), .ZN(_06109_ ) );
NAND3_X1 _13748_ ( .A1(_06107_ ), .A2(_05416_ ), .A3(\fc_addr [28] ), .ZN(_06110_ ) );
AOI21_X1 _13749_ ( .A(_06054_ ), .B1(_06109_ ), .B2(_06110_ ), .ZN(_06111_ ) );
AOI21_X2 _13750_ ( .A(_06111_ ), .B1(_05030_ ), .B2(_06055_ ), .ZN(_06112_ ) );
AOI211_X1 _13751_ ( .A(fanout_net_4 ), .B(_06098_ ), .C1(_06112_ ), .C2(_06069_ ), .ZN(_00522_ ) );
CLKBUF_X2 _13752_ ( .A(_00857_ ), .Z(_06113_ ) );
AND3_X1 _13753_ ( .A1(_01714_ ), .A2(_06113_ ), .A3(_01716_ ), .ZN(_06114_ ) );
AOI211_X1 _13754_ ( .A(_00770_ ), .B(_04722_ ), .C1(_04727_ ), .C2(_04769_ ), .ZN(_06115_ ) );
NAND3_X1 _13755_ ( .A1(_06081_ ), .A2(_06101_ ), .A3(_06104_ ), .ZN(_06116_ ) );
XNOR2_X1 _13756_ ( .A(_06116_ ), .B(\fc_addr [20] ), .ZN(_06117_ ) );
AOI21_X1 _13757_ ( .A(_06115_ ), .B1(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .B2(_06117_ ), .ZN(_06118_ ) );
AOI211_X1 _13758_ ( .A(fanout_net_4 ), .B(_06114_ ), .C1(_06118_ ), .C2(_06069_ ), .ZN(_00523_ ) );
AND3_X1 _13759_ ( .A1(_01773_ ), .A2(_06113_ ), .A3(_01775_ ), .ZN(_06119_ ) );
AOI211_X1 _13760_ ( .A(_00770_ ), .B(_04770_ ), .C1(_04798_ ), .C2(_04806_ ), .ZN(_06120_ ) );
NAND3_X1 _13761_ ( .A1(_06081_ ), .A2(\fc_addr [18] ), .A3(_06101_ ), .ZN(_06121_ ) );
XNOR2_X1 _13762_ ( .A(_06121_ ), .B(\fc_addr [19] ), .ZN(_06122_ ) );
AOI21_X1 _13763_ ( .A(_06120_ ), .B1(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .B2(_06122_ ), .ZN(_06123_ ) );
AOI211_X1 _13764_ ( .A(fanout_net_4 ), .B(_06119_ ), .C1(_06123_ ), .C2(_06069_ ), .ZN(_00524_ ) );
AOI211_X1 _13765_ ( .A(_00769_ ), .B(_04807_ ), .C1(_04834_ ), .C2(_04843_ ), .ZN(_06124_ ) );
XNOR2_X1 _13766_ ( .A(_06102_ ), .B(_05540_ ), .ZN(_06125_ ) );
AOI211_X1 _13767_ ( .A(_06113_ ), .B(_06124_ ), .C1(_00770_ ), .C2(_06125_ ), .ZN(_06126_ ) );
AOI211_X1 _13768_ ( .A(fanout_net_4 ), .B(_06126_ ), .C1(_00859_ ), .C2(_01842_ ), .ZN(_00525_ ) );
INV_X1 _13769_ ( .A(_06087_ ), .ZN(_06127_ ) );
OAI21_X1 _13770_ ( .A(_00769_ ), .B1(_06127_ ), .B2(_05657_ ), .ZN(_06128_ ) );
AOI21_X1 _13771_ ( .A(_06128_ ), .B1(_05657_ ), .B2(_06127_ ), .ZN(_06129_ ) );
BUF_X4 _13772_ ( .A(_06053_ ), .Z(_06130_ ) );
AOI211_X1 _13773_ ( .A(_06113_ ), .B(_06129_ ), .C1(_04880_ ), .C2(_06130_ ), .ZN(_06131_ ) );
AOI211_X1 _13774_ ( .A(fanout_net_4 ), .B(_06131_ ), .C1(_00859_ ), .C2(_01898_ ), .ZN(_00526_ ) );
AND3_X1 _13775_ ( .A1(_01948_ ), .A2(_06113_ ), .A3(_01949_ ), .ZN(_06132_ ) );
INV_X1 _13776_ ( .A(_06086_ ), .ZN(_06133_ ) );
OAI21_X1 _13777_ ( .A(_00770_ ), .B1(_06133_ ), .B2(_05439_ ), .ZN(_06134_ ) );
AOI21_X1 _13778_ ( .A(_06134_ ), .B1(_05439_ ), .B2(_06133_ ), .ZN(_06135_ ) );
AOI21_X1 _13779_ ( .A(_06135_ ), .B1(_04901_ ), .B2(_06055_ ), .ZN(_06136_ ) );
AOI211_X1 _13780_ ( .A(fanout_net_4 ), .B(_06132_ ), .C1(_06136_ ), .C2(_06069_ ), .ZN(_00527_ ) );
INV_X1 _13781_ ( .A(_06085_ ), .ZN(_06137_ ) );
OAI21_X1 _13782_ ( .A(_00769_ ), .B1(_06137_ ), .B2(_05661_ ), .ZN(_06138_ ) );
AOI21_X1 _13783_ ( .A(_06138_ ), .B1(_05661_ ), .B2(_06137_ ), .ZN(_06139_ ) );
AOI21_X1 _13784_ ( .A(_04902_ ), .B1(_04912_ ), .B2(_04935_ ), .ZN(_06140_ ) );
AOI211_X1 _13785_ ( .A(_06113_ ), .B(_06139_ ), .C1(_06140_ ), .C2(_06130_ ), .ZN(_06141_ ) );
AOI211_X1 _13786_ ( .A(fanout_net_4 ), .B(_06141_ ), .C1(_00859_ ), .C2(_01988_ ), .ZN(_00528_ ) );
INV_X1 _13787_ ( .A(_06084_ ), .ZN(_06142_ ) );
OAI21_X1 _13788_ ( .A(_00769_ ), .B1(_06142_ ), .B2(_05664_ ), .ZN(_06143_ ) );
AOI21_X1 _13789_ ( .A(_06143_ ), .B1(_05664_ ), .B2(_06142_ ), .ZN(_06144_ ) );
AOI21_X1 _13790_ ( .A(_04936_ ), .B1(_04939_ ), .B2(_04958_ ), .ZN(_06145_ ) );
AOI211_X1 _13791_ ( .A(_06113_ ), .B(_06144_ ), .C1(_06145_ ), .C2(_06130_ ), .ZN(_06146_ ) );
AOI211_X1 _13792_ ( .A(fanout_net_4 ), .B(_06146_ ), .C1(_00859_ ), .C2(_02044_ ), .ZN(_00529_ ) );
INV_X1 _13793_ ( .A(_06083_ ), .ZN(_06147_ ) );
OAI21_X1 _13794_ ( .A(_00769_ ), .B1(_06147_ ), .B2(_05425_ ), .ZN(_06148_ ) );
AOI21_X1 _13795_ ( .A(_06148_ ), .B1(_05425_ ), .B2(_06147_ ), .ZN(_06149_ ) );
AOI211_X1 _13796_ ( .A(_00857_ ), .B(_06149_ ), .C1(_04985_ ), .C2(_06130_ ), .ZN(_06150_ ) );
AOI211_X1 _13797_ ( .A(fanout_net_4 ), .B(_06150_ ), .C1(_00859_ ), .C2(_02091_ ), .ZN(_00530_ ) );
AND3_X1 _13798_ ( .A1(_02131_ ), .A2(_06113_ ), .A3(_02136_ ), .ZN(_06151_ ) );
INV_X1 _13799_ ( .A(_06081_ ), .ZN(_06152_ ) );
OAI21_X1 _13800_ ( .A(\fc_addr [12] ), .B1(_06152_ ), .B2(_06100_ ), .ZN(_06153_ ) );
NAND4_X1 _13801_ ( .A1(_06081_ ), .A2(_05516_ ), .A3(\fc_addr [11] ), .A4(\fc_addr [10] ), .ZN(_06154_ ) );
AOI21_X1 _13802_ ( .A(_06054_ ), .B1(_06153_ ), .B2(_06154_ ), .ZN(_06155_ ) );
AOI21_X1 _13803_ ( .A(_06155_ ), .B1(_05006_ ), .B2(_06055_ ), .ZN(_06156_ ) );
AOI211_X1 _13804_ ( .A(fanout_net_4 ), .B(_06151_ ), .C1(_06156_ ), .C2(_06069_ ), .ZN(_00531_ ) );
INV_X1 _13805_ ( .A(_06082_ ), .ZN(_06157_ ) );
OAI21_X1 _13806_ ( .A(_00769_ ), .B1(_06157_ ), .B2(_05533_ ), .ZN(_06158_ ) );
AOI21_X1 _13807_ ( .A(_06158_ ), .B1(_05533_ ), .B2(_06157_ ), .ZN(_06159_ ) );
AOI21_X1 _13808_ ( .A(_05031_ ), .B1(_05036_ ), .B2(_05055_ ), .ZN(_06160_ ) );
AOI211_X1 _13809_ ( .A(_00857_ ), .B(_06159_ ), .C1(_06160_ ), .C2(_06130_ ), .ZN(_06161_ ) );
AOI211_X1 _13810_ ( .A(fanout_net_4 ), .B(_06161_ ), .C1(_00859_ ), .C2(_02218_ ), .ZN(_00532_ ) );
OR2_X1 _13811_ ( .A1(_06107_ ), .A2(_05693_ ), .ZN(_06162_ ) );
NAND4_X1 _13812_ ( .A1(_06106_ ), .A2(_05693_ ), .A3(\fc_addr [27] ), .A4(\fc_addr [26] ), .ZN(_06163_ ) );
AOI21_X1 _13813_ ( .A(_06053_ ), .B1(_06162_ ), .B2(_06163_ ), .ZN(_06164_ ) );
AOI211_X1 _13814_ ( .A(_00857_ ), .B(_06164_ ), .C1(_05268_ ), .C2(_06130_ ), .ZN(_06165_ ) );
AOI211_X1 _13815_ ( .A(fanout_net_4 ), .B(_06165_ ), .C1(_00859_ ), .C2(_02716_ ), .ZN(_00533_ ) );
AND3_X1 _13816_ ( .A1(_02265_ ), .A2(_06113_ ), .A3(_02266_ ), .ZN(_06166_ ) );
OAI21_X1 _13817_ ( .A(_00770_ ), .B1(_06152_ ), .B2(_05676_ ), .ZN(_06167_ ) );
AOI21_X1 _13818_ ( .A(_06167_ ), .B1(_05676_ ), .B2(_06152_ ), .ZN(_06168_ ) );
AOI21_X1 _13819_ ( .A(_06168_ ), .B1(_05077_ ), .B2(_06055_ ), .ZN(_06169_ ) );
AOI211_X1 _13820_ ( .A(fanout_net_4 ), .B(_06166_ ), .C1(_06169_ ), .C2(_06069_ ), .ZN(_00534_ ) );
AND3_X1 _13821_ ( .A1(_02311_ ), .A2(_06113_ ), .A3(_02312_ ), .ZN(_06170_ ) );
INV_X1 _13822_ ( .A(_06080_ ), .ZN(_06171_ ) );
OAI21_X1 _13823_ ( .A(_00769_ ), .B1(_06171_ ), .B2(_05678_ ), .ZN(_06172_ ) );
AOI21_X1 _13824_ ( .A(_06172_ ), .B1(_05678_ ), .B2(_06171_ ), .ZN(_06173_ ) );
AOI21_X1 _13825_ ( .A(_05078_ ), .B1(_05084_ ), .B2(_05103_ ), .ZN(_06174_ ) );
AOI21_X1 _13826_ ( .A(_06173_ ), .B1(_06174_ ), .B2(_06055_ ), .ZN(_06175_ ) );
AOI211_X1 _13827_ ( .A(fanout_net_4 ), .B(_06170_ ), .C1(_06175_ ), .C2(_06069_ ), .ZN(_00535_ ) );
AOI21_X1 _13828_ ( .A(\fc_addr [8] ), .B1(_06078_ ), .B2(\fc_addr [7] ), .ZN(_06176_ ) );
NOR3_X1 _13829_ ( .A1(_06080_ ), .A2(_06054_ ), .A3(_06176_ ), .ZN(_06177_ ) );
AOI21_X1 _13830_ ( .A(_06177_ ), .B1(_05120_ ), .B2(_06055_ ), .ZN(_06178_ ) );
NAND2_X1 _13831_ ( .A1(_00857_ ), .A2(_00771_ ), .ZN(_06179_ ) );
BUF_X4 _13832_ ( .A(_06179_ ), .Z(_06180_ ) );
OAI22_X1 _13833_ ( .A1(_06178_ ), .A2(_04455_ ), .B1(_02354_ ), .B2(_06180_ ), .ZN(_00536_ ) );
XNOR2_X1 _13834_ ( .A(_06078_ ), .B(\fc_addr [7] ), .ZN(_06181_ ) );
MUX2_X1 _13835_ ( .A(_06181_ ), .B(_05145_ ), .S(_06054_ ), .Z(_06182_ ) );
OAI22_X1 _13836_ ( .A1(_06182_ ), .A2(_04455_ ), .B1(_02398_ ), .B2(_06180_ ), .ZN(_00537_ ) );
AND2_X1 _13837_ ( .A1(_02447_ ), .A2(_02448_ ), .ZN(_06183_ ) );
NOR2_X1 _13838_ ( .A1(_06077_ ), .A2(\fc_addr [6] ), .ZN(_06184_ ) );
NOR3_X1 _13839_ ( .A1(_06078_ ), .A2(_06184_ ), .A3(_06053_ ), .ZN(_06185_ ) );
AOI21_X1 _13840_ ( .A(_06185_ ), .B1(_05166_ ), .B2(_06055_ ), .ZN(_06186_ ) );
OAI22_X1 _13841_ ( .A1(_06183_ ), .A2(_06180_ ), .B1(_06186_ ), .B2(_00880_ ), .ZN(_00538_ ) );
INV_X1 _13842_ ( .A(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B ), .ZN(_06187_ ) );
AOI21_X1 _13843_ ( .A(\fc_addr [5] ), .B1(_05731_ ), .B2(_06187_ ), .ZN(_06188_ ) );
AND4_X1 _13844_ ( .A1(\fc_addr [5] ), .A2(_06187_ ), .A3(\fc_addr [3] ), .A4(\fc_addr [2] ), .ZN(_06189_ ) );
NOR3_X1 _13845_ ( .A1(_06188_ ), .A2(_06054_ ), .A3(_06189_ ), .ZN(_06190_ ) );
AOI21_X1 _13846_ ( .A(_06190_ ), .B1(_05187_ ), .B2(_06055_ ), .ZN(_06191_ ) );
OAI22_X1 _13847_ ( .A1(_06191_ ), .A2(_04455_ ), .B1(_04459_ ), .B2(_06180_ ), .ZN(_00539_ ) );
XNOR2_X1 _13848_ ( .A(_05729_ ), .B(\fc_addr [4] ), .ZN(_06192_ ) );
NAND2_X1 _13849_ ( .A1(_06192_ ), .A2(_00769_ ), .ZN(_06193_ ) );
OAI21_X1 _13850_ ( .A(_06193_ ), .B1(_05204_ ), .B2(_00770_ ), .ZN(_06194_ ) );
MUX2_X1 _13851_ ( .A(_06194_ ), .B(_02558_ ), .S(_00857_ ), .Z(_06195_ ) );
NOR2_X1 _13852_ ( .A1(_06195_ ), .A2(reset ), .ZN(_00540_ ) );
XNOR2_X1 _13853_ ( .A(\fc_addr [3] ), .B(\fc_addr [2] ), .ZN(_06196_ ) );
MUX2_X1 _13854_ ( .A(_06196_ ), .B(_05228_ ), .S(_06054_ ), .Z(_06197_ ) );
AND2_X1 _13855_ ( .A1(_02609_ ), .A2(_02610_ ), .ZN(_06198_ ) );
OAI22_X1 _13856_ ( .A1(_06197_ ), .A2(_04455_ ), .B1(_06198_ ), .B2(_06180_ ), .ZN(_00541_ ) );
OAI21_X1 _13857_ ( .A(_00772_ ), .B1(_00000_ ), .B2(\fc_addr [4] ), .ZN(_06199_ ) );
AOI21_X1 _13858_ ( .A(_06199_ ), .B1(_06195_ ), .B2(_00000_ ), .ZN(_00542_ ) );
OR2_X1 _13859_ ( .A1(_06054_ ), .A2(\u_ifu.pc_$_SDFFE_PP0N__Q_28_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06200_ ) );
OAI211_X1 _13860_ ( .A(_00878_ ), .B(_06200_ ), .C1(_05242_ ), .C2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06201_ ) );
OAI21_X1 _13861_ ( .A(_06201_ ), .B1(_02675_ ), .B2(_06180_ ), .ZN(_00543_ ) );
NAND3_X1 _13862_ ( .A1(_06102_ ), .A2(\fc_addr [26] ), .A3(_06105_ ), .ZN(_06202_ ) );
NAND2_X1 _13863_ ( .A1(_06202_ ), .A2(\fc_addr [27] ), .ZN(_06203_ ) );
NAND4_X1 _13864_ ( .A1(_06102_ ), .A2(_05462_ ), .A3(\fc_addr [26] ), .A4(_06105_ ), .ZN(_06204_ ) );
NAND3_X1 _13865_ ( .A1(_06203_ ), .A2(_00770_ ), .A3(_06204_ ), .ZN(_06205_ ) );
OAI211_X1 _13866_ ( .A(_00878_ ), .B(_06205_ ), .C1(_05312_ ), .C2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06206_ ) );
AND2_X1 _13867_ ( .A1(_02859_ ), .A2(_02860_ ), .ZN(_06207_ ) );
OAI21_X1 _13868_ ( .A(_06206_ ), .B1(_06207_ ), .B2(_06180_ ), .ZN(_00544_ ) );
OAI21_X1 _13869_ ( .A(_00878_ ), .B1(_05330_ ), .B2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06208_ ) );
AOI21_X1 _13870_ ( .A(_05469_ ), .B1(_06102_ ), .B2(_06105_ ), .ZN(_06209_ ) );
AND4_X1 _13871_ ( .A1(_05469_ ), .A2(_06081_ ), .A3(_06101_ ), .A4(_06105_ ), .ZN(_06210_ ) );
NOR3_X1 _13872_ ( .A1(_06209_ ), .A2(_06130_ ), .A3(_06210_ ), .ZN(_06211_ ) );
OAI22_X1 _13873_ ( .A1(_06208_ ), .A2(_06211_ ), .B1(_02898_ ), .B2(_06179_ ), .ZN(_00545_ ) );
AOI211_X1 _13874_ ( .A(_00770_ ), .B(_05331_ ), .C1(_05334_ ), .C2(_05346_ ), .ZN(_06212_ ) );
AND3_X1 _13875_ ( .A1(_06104_ ), .A2(\fc_addr [21] ), .A3(\fc_addr [20] ), .ZN(_06213_ ) );
AND2_X1 _13876_ ( .A1(_06102_ ), .A2(_06213_ ), .ZN(_06214_ ) );
AND3_X1 _13877_ ( .A1(_06214_ ), .A2(\fc_addr [23] ), .A3(\fc_addr [22] ), .ZN(_06215_ ) );
NAND2_X1 _13878_ ( .A1(_06215_ ), .A2(\fc_addr [24] ), .ZN(_06216_ ) );
NAND2_X1 _13879_ ( .A1(_06216_ ), .A2(\fc_addr [25] ), .ZN(_06217_ ) );
NAND3_X1 _13880_ ( .A1(_06215_ ), .A2(_05458_ ), .A3(\fc_addr [24] ), .ZN(_06218_ ) );
AOI21_X1 _13881_ ( .A(_06054_ ), .B1(_06217_ ), .B2(_06218_ ), .ZN(_06219_ ) );
OAI211_X1 _13882_ ( .A(_00772_ ), .B(_06068_ ), .C1(_06212_ ), .C2(_06219_ ), .ZN(_06220_ ) );
AND2_X1 _13883_ ( .A1(_02933_ ), .A2(_02934_ ), .ZN(_06221_ ) );
OAI21_X1 _13884_ ( .A(_06220_ ), .B1(_06221_ ), .B2(_06180_ ), .ZN(_00546_ ) );
OAI21_X1 _13885_ ( .A(_00878_ ), .B1(_05363_ ), .B2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06222_ ) );
NOR2_X1 _13886_ ( .A1(_06215_ ), .A2(_05708_ ), .ZN(_06223_ ) );
AND4_X1 _13887_ ( .A1(_05708_ ), .A2(_06214_ ), .A3(\fc_addr [23] ), .A4(\fc_addr [22] ), .ZN(_06224_ ) );
NOR3_X1 _13888_ ( .A1(_06223_ ), .A2(_06130_ ), .A3(_06224_ ), .ZN(_06225_ ) );
AND2_X1 _13889_ ( .A1(_02977_ ), .A2(_02978_ ), .ZN(_06226_ ) );
OAI22_X1 _13890_ ( .A1(_06222_ ), .A2(_06225_ ), .B1(_06226_ ), .B2(_06179_ ), .ZN(_00547_ ) );
NAND3_X1 _13891_ ( .A1(_06102_ ), .A2(\fc_addr [22] ), .A3(_06213_ ), .ZN(_06227_ ) );
XNOR2_X1 _13892_ ( .A(_06227_ ), .B(\fc_addr [23] ), .ZN(_06228_ ) );
OR2_X1 _13893_ ( .A1(_06228_ ), .A2(_06053_ ), .ZN(_06229_ ) );
OAI211_X2 _13894_ ( .A(_00878_ ), .B(_06229_ ), .C1(_05382_ ), .C2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06230_ ) );
OAI21_X1 _13895_ ( .A(_06230_ ), .B1(_03024_ ), .B2(_06180_ ), .ZN(_00548_ ) );
XNOR2_X1 _13896_ ( .A(_06214_ ), .B(_05451_ ), .ZN(_06231_ ) );
MUX2_X1 _13897_ ( .A(_06231_ ), .B(_05399_ ), .S(_06053_ ), .Z(_06232_ ) );
AND3_X1 _13898_ ( .A1(_06232_ ), .A2(_00772_ ), .A3(_06068_ ), .ZN(_06233_ ) );
AOI21_X1 _13899_ ( .A(_06179_ ), .B1(_03069_ ), .B2(_03070_ ), .ZN(_06234_ ) );
OR2_X1 _13900_ ( .A1(_06233_ ), .A2(_06234_ ), .ZN(_00549_ ) );
NOR2_X1 _13901_ ( .A1(_06116_ ), .A2(_05530_ ), .ZN(_06235_ ) );
XNOR2_X1 _13902_ ( .A(_06235_ ), .B(_05650_ ), .ZN(_06236_ ) );
MUX2_X2 _13903_ ( .A(_06236_ ), .B(_04721_ ), .S(_06053_ ), .Z(_06237_ ) );
AND3_X2 _13904_ ( .A1(_06237_ ), .A2(_00771_ ), .A3(_06068_ ), .ZN(_06238_ ) );
AOI21_X1 _13905_ ( .A(_06179_ ), .B1(_01658_ ), .B2(_01659_ ), .ZN(_06239_ ) );
OR2_X2 _13906_ ( .A1(_06238_ ), .A2(_06239_ ), .ZN(_00550_ ) );
NAND3_X1 _13907_ ( .A1(_00865_ ), .A2(_00771_ ), .A3(_06053_ ), .ZN(_06240_ ) );
OR3_X1 _13908_ ( .A1(_05288_ ), .A2(_05289_ ), .A3(_06240_ ), .ZN(_06241_ ) );
OAI21_X1 _13909_ ( .A(_06241_ ), .B1(_02767_ ), .B2(_06180_ ), .ZN(_00551_ ) );
OAI22_X1 _13910_ ( .A1(_04210_ ), .A2(_06240_ ), .B1(_02822_ ), .B2(_06179_ ), .ZN(_00552_ ) );
AND2_X1 _13911_ ( .A1(_01470_ ), .A2(_01473_ ), .ZN(_06242_ ) );
OAI21_X1 _13912_ ( .A(_06068_ ), .B1(_04592_ ), .B2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(_06243_ ) );
AND2_X1 _13913_ ( .A1(_06094_ ), .A2(\fc_addr [28] ), .ZN(_06244_ ) );
NAND4_X1 _13914_ ( .A1(_06244_ ), .A2(\fc_addr [31] ), .A3(\fc_addr [30] ), .A4(\fc_addr [29] ), .ZN(_06245_ ) );
OAI21_X1 _13915_ ( .A(_05442_ ), .B1(_06095_ ), .B2(_05525_ ), .ZN(_06246_ ) );
AOI21_X1 _13916_ ( .A(_06130_ ), .B1(_06245_ ), .B2(_06246_ ), .ZN(_06247_ ) );
OAI221_X1 _13917_ ( .A(_00773_ ), .B1(_06069_ ), .B2(_06242_ ), .C1(_06243_ ), .C2(_06247_ ), .ZN(_00553_ ) );
OR2_X1 _13918_ ( .A1(_01280_ ), .A2(\u_lsu.reading ), .ZN(_06248_ ) );
NOR4_X1 _13919_ ( .A1(_06066_ ), .A2(reset ), .A3(_06067_ ), .A4(_06248_ ), .ZN(_00554_ ) );
OAI21_X1 _13920_ ( .A(\u_arbiter.wvalid ), .B1(_01170_ ), .B2(\u_arbiter.working ), .ZN(_06249_ ) );
NOR4_X1 _13921_ ( .A1(flush_$_OR__Y_B ), .A2(\u_lsu.writing ), .A3(_05717_ ), .A4(_06249_ ), .ZN(_00555_ ) );
AND2_X1 _13922_ ( .A1(\u_lsu.rcount [0] ), .A2(\u_lsu.rcount [1] ), .ZN(_06250_ ) );
AND2_X1 _13923_ ( .A1(_06250_ ), .A2(\u_lsu.rcount [2] ), .ZN(_06251_ ) );
AND2_X1 _13924_ ( .A1(_06251_ ), .A2(\u_lsu.rcount [3] ), .ZN(_06252_ ) );
AND2_X1 _13925_ ( .A1(_06252_ ), .A2(\u_lsu.rcount [4] ), .ZN(_06253_ ) );
AND2_X1 _13926_ ( .A1(_06253_ ), .A2(\u_lsu.rcount [5] ), .ZN(_06254_ ) );
AND2_X1 _13927_ ( .A1(_06254_ ), .A2(\u_lsu.rcount [6] ), .ZN(_06255_ ) );
XNOR2_X1 _13928_ ( .A(_06255_ ), .B(\u_lsu.rcount [7] ), .ZN(_06256_ ) );
NOR2_X1 _13929_ ( .A1(_04461_ ), .A2(_06256_ ), .ZN(_00556_ ) );
OAI211_X1 _13930_ ( .A(_04454_ ), .B(_06061_ ), .C1(\u_lsu.rcount [6] ), .C2(_06254_ ), .ZN(_06257_ ) );
NOR2_X1 _13931_ ( .A1(_06257_ ), .A2(_06255_ ), .ZN(_00557_ ) );
OAI211_X1 _13932_ ( .A(_04454_ ), .B(_06061_ ), .C1(\u_lsu.rcount [5] ), .C2(_06253_ ), .ZN(_06258_ ) );
NOR2_X1 _13933_ ( .A1(_06258_ ), .A2(_06254_ ), .ZN(_00558_ ) );
OAI211_X1 _13934_ ( .A(_04454_ ), .B(_06061_ ), .C1(\u_lsu.rcount [4] ), .C2(_06252_ ), .ZN(_06259_ ) );
NOR2_X1 _13935_ ( .A1(_06259_ ), .A2(_06253_ ), .ZN(_00559_ ) );
OAI211_X1 _13936_ ( .A(_04454_ ), .B(_06068_ ), .C1(\u_lsu.rcount [3] ), .C2(_06251_ ), .ZN(_06260_ ) );
NOR2_X1 _13937_ ( .A1(_06260_ ), .A2(_06252_ ), .ZN(_00560_ ) );
OAI211_X1 _13938_ ( .A(_04454_ ), .B(_06068_ ), .C1(\u_lsu.rcount [2] ), .C2(_06250_ ), .ZN(_06261_ ) );
NOR2_X1 _13939_ ( .A1(_06261_ ), .A2(_06251_ ), .ZN(_00561_ ) );
NOR2_X1 _13940_ ( .A1(\u_lsu.rcount [0] ), .A2(\u_lsu.rcount [1] ), .ZN(_06262_ ) );
NOR4_X1 _13941_ ( .A1(flush_$_OR__Y_B ), .A2(_00882_ ), .A3(_06250_ ), .A4(_06262_ ), .ZN(_00562_ ) );
NOR4_X1 _13942_ ( .A1(\u_lsu.rcount [6] ), .A2(\u_lsu.rcount [5] ), .A3(\u_lsu.rcount [4] ), .A4(\u_lsu.rcount [7] ), .ZN(_06263_ ) );
NOR4_X1 _13943_ ( .A1(\u_lsu.rcount [3] ), .A2(\u_lsu.rcount [2] ), .A3(\u_lsu.rcount [0] ), .A4(\u_lsu.rcount [1] ), .ZN(_06264_ ) );
AND2_X1 _13944_ ( .A1(_06263_ ), .A2(_06264_ ), .ZN(_06265_ ) );
NOR4_X1 _13945_ ( .A1(flush_$_OR__Y_B ), .A2(\u_lsu.rcount [0] ), .A3(_05717_ ), .A4(_06265_ ), .ZN(_00563_ ) );
NAND3_X4 _13946_ ( .A1(\u_lsu.u_clint.mtime [1] ), .A2(\u_lsu.u_clint.mtime [2] ), .A3(\u_lsu.u_clint.mtime [0] ), .ZN(_06266_ ) );
NOR2_X4 _13947_ ( .A1(_06266_ ), .A2(_02577_ ), .ZN(_06267_ ) );
AND2_X4 _13948_ ( .A1(\u_lsu.u_clint.mtime [5] ), .A2(\u_lsu.u_clint.mtime [4] ), .ZN(_06268_ ) );
AND2_X4 _13949_ ( .A1(_06267_ ), .A2(_06268_ ), .ZN(_06269_ ) );
INV_X4 _13950_ ( .A(_06269_ ), .ZN(_06270_ ) );
NAND2_X4 _13951_ ( .A1(\u_lsu.u_clint.mtime [7] ), .A2(\u_lsu.u_clint.mtime [6] ), .ZN(_06271_ ) );
NOR2_X4 _13952_ ( .A1(_06270_ ), .A2(_06271_ ), .ZN(_06272_ ) );
AND2_X2 _13953_ ( .A1(\u_lsu.u_clint.mtime [9] ), .A2(\u_lsu.u_clint.mtime [8] ), .ZN(_06273_ ) );
AND3_X4 _13954_ ( .A1(_06272_ ), .A2(\u_lsu.u_clint.mtime [10] ), .A3(_06273_ ), .ZN(_06274_ ) );
AND3_X4 _13955_ ( .A1(_06274_ ), .A2(\u_lsu.u_clint.mtime [11] ), .A3(\u_lsu.u_clint.mtime [12] ), .ZN(_06275_ ) );
AND2_X4 _13956_ ( .A1(_06275_ ), .A2(\u_lsu.u_clint.mtime [13] ), .ZN(_06276_ ) );
AND2_X1 _13957_ ( .A1(\u_lsu.u_clint.mtime [15] ), .A2(\u_lsu.u_clint.mtime [14] ), .ZN(_06277_ ) );
AND2_X4 _13958_ ( .A1(_06276_ ), .A2(_06277_ ), .ZN(_06278_ ) );
AND2_X1 _13959_ ( .A1(\u_lsu.u_clint.mtime [17] ), .A2(\u_lsu.u_clint.mtime [16] ), .ZN(_06279_ ) );
AND2_X4 _13960_ ( .A1(_06278_ ), .A2(_06279_ ), .ZN(_06280_ ) );
AND2_X1 _13961_ ( .A1(\u_lsu.u_clint.mtime [19] ), .A2(\u_lsu.u_clint.mtime [18] ), .ZN(_06281_ ) );
AND2_X4 _13962_ ( .A1(_06280_ ), .A2(_06281_ ), .ZN(_06282_ ) );
AND2_X1 _13963_ ( .A1(\u_lsu.u_clint.mtime [21] ), .A2(\u_lsu.u_clint.mtime [20] ), .ZN(_06283_ ) );
AND2_X4 _13964_ ( .A1(_06282_ ), .A2(_06283_ ), .ZN(_06284_ ) );
AND2_X1 _13965_ ( .A1(\u_lsu.u_clint.mtime [23] ), .A2(\u_lsu.u_clint.mtime [22] ), .ZN(_06285_ ) );
AND2_X4 _13966_ ( .A1(_06284_ ), .A2(_06285_ ), .ZN(_06286_ ) );
AND2_X1 _13967_ ( .A1(\u_lsu.u_clint.mtime [25] ), .A2(\u_lsu.u_clint.mtime [24] ), .ZN(_06287_ ) );
AND2_X4 _13968_ ( .A1(_06286_ ), .A2(_06287_ ), .ZN(_06288_ ) );
AND2_X1 _13969_ ( .A1(\u_lsu.u_clint.mtime [27] ), .A2(\u_lsu.u_clint.mtime [26] ), .ZN(_06289_ ) );
AND2_X4 _13970_ ( .A1(_06288_ ), .A2(_06289_ ), .ZN(_06290_ ) );
AND2_X1 _13971_ ( .A1(\u_lsu.u_clint.mtime [29] ), .A2(\u_lsu.u_clint.mtime [28] ), .ZN(_06291_ ) );
AND2_X4 _13972_ ( .A1(_06290_ ), .A2(_06291_ ), .ZN(_06292_ ) );
AND2_X1 _13973_ ( .A1(\u_lsu.u_clint.mtime [31] ), .A2(\u_lsu.u_clint.mtime [30] ), .ZN(_06293_ ) );
AND2_X4 _13974_ ( .A1(_06292_ ), .A2(_06293_ ), .ZN(_06294_ ) );
AND2_X1 _13975_ ( .A1(\u_lsu.u_clint.mtime [33] ), .A2(\u_lsu.u_clint.mtime [32] ), .ZN(_06295_ ) );
AND2_X4 _13976_ ( .A1(_06294_ ), .A2(_06295_ ), .ZN(_06296_ ) );
AND2_X1 _13977_ ( .A1(\u_lsu.u_clint.mtime [35] ), .A2(\u_lsu.u_clint.mtime [34] ), .ZN(_06297_ ) );
AND2_X4 _13978_ ( .A1(_06296_ ), .A2(_06297_ ), .ZN(_06298_ ) );
AND2_X1 _13979_ ( .A1(\u_lsu.u_clint.mtime [37] ), .A2(\u_lsu.u_clint.mtime [36] ), .ZN(_06299_ ) );
AND3_X1 _13980_ ( .A1(_06299_ ), .A2(\u_lsu.u_clint.mtime [39] ), .A3(\u_lsu.u_clint.mtime [38] ), .ZN(_06300_ ) );
AND2_X4 _13981_ ( .A1(_06298_ ), .A2(_06300_ ), .ZN(_06301_ ) );
AND2_X1 _13982_ ( .A1(\u_lsu.u_clint.mtime [41] ), .A2(\u_lsu.u_clint.mtime [40] ), .ZN(_06302_ ) );
AND2_X4 _13983_ ( .A1(_06301_ ), .A2(_06302_ ), .ZN(_06303_ ) );
AND2_X1 _13984_ ( .A1(\u_lsu.u_clint.mtime [43] ), .A2(\u_lsu.u_clint.mtime [42] ), .ZN(_06304_ ) );
AND2_X4 _13985_ ( .A1(_06303_ ), .A2(_06304_ ), .ZN(_06305_ ) );
AND2_X1 _13986_ ( .A1(\u_lsu.u_clint.mtime [45] ), .A2(\u_lsu.u_clint.mtime [44] ), .ZN(_06306_ ) );
AND3_X1 _13987_ ( .A1(_06306_ ), .A2(\u_lsu.u_clint.mtime [47] ), .A3(\u_lsu.u_clint.mtime [46] ), .ZN(_06307_ ) );
AND2_X4 _13988_ ( .A1(_06305_ ), .A2(_06307_ ), .ZN(_06308_ ) );
AND2_X1 _13989_ ( .A1(\u_lsu.u_clint.mtime [49] ), .A2(\u_lsu.u_clint.mtime [48] ), .ZN(_06309_ ) );
AND2_X4 _13990_ ( .A1(_06308_ ), .A2(_06309_ ), .ZN(_06310_ ) );
AND2_X1 _13991_ ( .A1(\u_lsu.u_clint.mtime [51] ), .A2(\u_lsu.u_clint.mtime [50] ), .ZN(_06311_ ) );
AND2_X4 _13992_ ( .A1(_06310_ ), .A2(_06311_ ), .ZN(_06312_ ) );
AND2_X1 _13993_ ( .A1(\u_lsu.u_clint.mtime [53] ), .A2(\u_lsu.u_clint.mtime [52] ), .ZN(_06313_ ) );
AND2_X4 _13994_ ( .A1(_06312_ ), .A2(_06313_ ), .ZN(_06314_ ) );
AND2_X1 _13995_ ( .A1(\u_lsu.u_clint.mtime [55] ), .A2(\u_lsu.u_clint.mtime [54] ), .ZN(_06315_ ) );
AND2_X4 _13996_ ( .A1(_06314_ ), .A2(_06315_ ), .ZN(_06316_ ) );
AND2_X1 _13997_ ( .A1(\u_lsu.u_clint.mtime [57] ), .A2(\u_lsu.u_clint.mtime [56] ), .ZN(_06317_ ) );
AND2_X4 _13998_ ( .A1(_06316_ ), .A2(_06317_ ), .ZN(_06318_ ) );
AND2_X1 _13999_ ( .A1(\u_lsu.u_clint.mtime [59] ), .A2(\u_lsu.u_clint.mtime [58] ), .ZN(_06319_ ) );
AND2_X4 _14000_ ( .A1(_06318_ ), .A2(_06319_ ), .ZN(_06320_ ) );
NAND3_X4 _14001_ ( .A1(_06320_ ), .A2(\u_lsu.u_clint.mtime [61] ), .A3(\u_lsu.u_clint.mtime [60] ), .ZN(_06321_ ) );
NOR2_X4 _14002_ ( .A1(_06321_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ), .ZN(_06322_ ) );
AND2_X2 _14003_ ( .A1(_06322_ ), .A2(\u_lsu.u_clint.mtime [63] ), .ZN(_06323_ ) );
OAI21_X1 _14004_ ( .A(_04476_ ), .B1(_06322_ ), .B2(\u_lsu.u_clint.mtime [63] ), .ZN(_06324_ ) );
NOR2_X1 _14005_ ( .A1(_06323_ ), .A2(_06324_ ), .ZN(_00564_ ) );
INV_X1 _14006_ ( .A(_06272_ ), .ZN(_06325_ ) );
AND3_X1 _14007_ ( .A1(_06273_ ), .A2(\u_lsu.u_clint.mtime [11] ), .A3(\u_lsu.u_clint.mtime [10] ), .ZN(_06326_ ) );
NAND4_X1 _14008_ ( .A1(_06326_ ), .A2(\u_lsu.u_clint.mtime [13] ), .A3(\u_lsu.u_clint.mtime [12] ), .A4(_06277_ ), .ZN(_06327_ ) );
NOR2_X1 _14009_ ( .A1(_06325_ ), .A2(_06327_ ), .ZN(_06328_ ) );
AND2_X1 _14010_ ( .A1(_06281_ ), .A2(_06279_ ), .ZN(_06329_ ) );
AND3_X1 _14011_ ( .A1(_06329_ ), .A2(_06285_ ), .A3(_06283_ ), .ZN(_06330_ ) );
AND2_X1 _14012_ ( .A1(_06289_ ), .A2(_06287_ ), .ZN(_06331_ ) );
AND4_X1 _14013_ ( .A1(_06293_ ), .A2(_06330_ ), .A3(_06291_ ), .A4(_06331_ ), .ZN(_06332_ ) );
AND2_X1 _14014_ ( .A1(_06328_ ), .A2(_06332_ ), .ZN(_06333_ ) );
AND2_X1 _14015_ ( .A1(_06304_ ), .A2(_06302_ ), .ZN(_06334_ ) );
AND2_X1 _14016_ ( .A1(_06297_ ), .A2(_06295_ ), .ZN(_06335_ ) );
AND4_X1 _14017_ ( .A1(_06307_ ), .A2(_06300_ ), .A3(_06334_ ), .A4(_06335_ ), .ZN(_06336_ ) );
AND2_X1 _14018_ ( .A1(_06333_ ), .A2(_06336_ ), .ZN(_06337_ ) );
AND4_X1 _14019_ ( .A1(_06315_ ), .A2(_06313_ ), .A3(_06311_ ), .A4(_06309_ ), .ZN(_06338_ ) );
AND2_X1 _14020_ ( .A1(_06337_ ), .A2(_06338_ ), .ZN(_06339_ ) );
AND4_X1 _14021_ ( .A1(\u_lsu.u_clint.mtime [59] ), .A2(\u_lsu.u_clint.mtime [57] ), .A3(\u_lsu.u_clint.mtime [58] ), .A4(\u_lsu.u_clint.mtime [56] ), .ZN(_06340_ ) );
AND2_X1 _14022_ ( .A1(_06339_ ), .A2(_06340_ ), .ZN(_06341_ ) );
AND3_X1 _14023_ ( .A1(_06341_ ), .A2(\u_lsu.u_clint.mtime [61] ), .A3(\u_lsu.u_clint.mtime [60] ), .ZN(_06342_ ) );
XNOR2_X1 _14024_ ( .A(_06342_ ), .B(\u_lsu.u_clint.mtime [62] ), .ZN(_06343_ ) );
NOR2_X1 _14025_ ( .A1(_06343_ ), .A2(_04472_ ), .ZN(_00565_ ) );
AND3_X1 _14026_ ( .A1(_06310_ ), .A2(_01680_ ), .A3(_06311_ ), .ZN(_06344_ ) );
OAI21_X1 _14027_ ( .A(_05622_ ), .B1(_06344_ ), .B2(\u_lsu.u_clint.mtime [53] ), .ZN(_06345_ ) );
AND4_X1 _14028_ ( .A1(\u_lsu.u_clint.mtime [53] ), .A2(_06310_ ), .A3(_01680_ ), .A4(_06311_ ), .ZN(_06346_ ) );
NOR2_X1 _14029_ ( .A1(_06345_ ), .A2(_06346_ ), .ZN(_00566_ ) );
AND2_X1 _14030_ ( .A1(_06311_ ), .A2(_06309_ ), .ZN(_06347_ ) );
AND2_X1 _14031_ ( .A1(_06337_ ), .A2(_06347_ ), .ZN(_06348_ ) );
XNOR2_X1 _14032_ ( .A(_06348_ ), .B(\u_lsu.u_clint.mtime [52] ), .ZN(_06349_ ) );
NOR2_X1 _14033_ ( .A1(_06349_ ), .A2(_04472_ ), .ZN(_00567_ ) );
INV_X1 _14034_ ( .A(_06310_ ), .ZN(_06350_ ) );
NOR2_X1 _14035_ ( .A1(_06350_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ), .ZN(_06351_ ) );
AND2_X1 _14036_ ( .A1(_06351_ ), .A2(\u_lsu.u_clint.mtime [51] ), .ZN(_06352_ ) );
OAI21_X1 _14037_ ( .A(_04476_ ), .B1(_06351_ ), .B2(\u_lsu.u_clint.mtime [51] ), .ZN(_06353_ ) );
NOR2_X1 _14038_ ( .A1(_06352_ ), .A2(_06353_ ), .ZN(_00568_ ) );
AND3_X1 _14039_ ( .A1(_06333_ ), .A2(_06309_ ), .A3(_06336_ ), .ZN(_06354_ ) );
XNOR2_X1 _14040_ ( .A(_06354_ ), .B(\u_lsu.u_clint.mtime [50] ), .ZN(_06355_ ) );
NOR2_X1 _14041_ ( .A1(_06355_ ), .A2(_04472_ ), .ZN(_00569_ ) );
AND3_X1 _14042_ ( .A1(_06305_ ), .A2(_01916_ ), .A3(_06307_ ), .ZN(_06356_ ) );
OAI21_X1 _14043_ ( .A(_05622_ ), .B1(_06356_ ), .B2(\u_lsu.u_clint.mtime [49] ), .ZN(_06357_ ) );
AND4_X1 _14044_ ( .A1(\u_lsu.u_clint.mtime [49] ), .A2(_06305_ ), .A3(_01916_ ), .A4(_06307_ ), .ZN(_06358_ ) );
NOR2_X1 _14045_ ( .A1(_06357_ ), .A2(_06358_ ), .ZN(_00570_ ) );
INV_X1 _14046_ ( .A(_06328_ ), .ZN(_06359_ ) );
INV_X1 _14047_ ( .A(_06332_ ), .ZN(_06360_ ) );
INV_X1 _14048_ ( .A(_06336_ ), .ZN(_06361_ ) );
OR4_X1 _14049_ ( .A1(\u_lsu.u_clint.mtime [48] ), .A2(_06359_ ), .A3(_06360_ ), .A4(_06361_ ), .ZN(_06362_ ) );
INV_X1 _14050_ ( .A(_06333_ ), .ZN(_06363_ ) );
OAI21_X1 _14051_ ( .A(\u_lsu.u_clint.mtime [48] ), .B1(_06363_ ), .B2(_06361_ ), .ZN(_06364_ ) );
AOI21_X1 _14052_ ( .A(_04462_ ), .B1(_06362_ ), .B2(_06364_ ), .ZN(_00571_ ) );
NAND3_X1 _14053_ ( .A1(_06303_ ), .A2(\u_lsu.u_clint.mtime [44] ), .A3(_06304_ ), .ZN(_06365_ ) );
NOR3_X1 _14054_ ( .A1(_06365_ ), .A2(_02056_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ), .ZN(_06366_ ) );
OAI21_X1 _14055_ ( .A(_05622_ ), .B1(_06366_ ), .B2(\u_lsu.u_clint.mtime [47] ), .ZN(_06367_ ) );
NOR4_X1 _14056_ ( .A1(_06365_ ), .A2(_01230_ ), .A3(_02056_ ), .A4(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ), .ZN(_06368_ ) );
NOR2_X1 _14057_ ( .A1(_06367_ ), .A2(_06368_ ), .ZN(_00572_ ) );
AND2_X1 _14058_ ( .A1(_06300_ ), .A2(_06335_ ), .ZN(_06369_ ) );
AND2_X1 _14059_ ( .A1(_06333_ ), .A2(_06369_ ), .ZN(_06370_ ) );
AND3_X1 _14060_ ( .A1(_06370_ ), .A2(_06306_ ), .A3(_06334_ ), .ZN(_06371_ ) );
XNOR2_X1 _14061_ ( .A(_06371_ ), .B(\u_lsu.u_clint.mtime [46] ), .ZN(_06372_ ) );
BUF_X4 _14062_ ( .A(_02455_ ), .Z(_06373_ ) );
NOR2_X1 _14063_ ( .A1(_06372_ ), .A2(_06373_ ), .ZN(_00573_ ) );
NAND3_X1 _14064_ ( .A1(_06303_ ), .A2(_02102_ ), .A3(_06304_ ), .ZN(_06374_ ) );
AOI21_X1 _14065_ ( .A(_02455_ ), .B1(_06374_ ), .B2(_02056_ ), .ZN(_06375_ ) );
NAND4_X1 _14066_ ( .A1(_06303_ ), .A2(\u_lsu.u_clint.mtime [45] ), .A3(_02102_ ), .A4(_06304_ ), .ZN(_06376_ ) );
AND2_X1 _14067_ ( .A1(_06375_ ), .A2(_06376_ ), .ZN(_00574_ ) );
AND2_X1 _14068_ ( .A1(_06370_ ), .A2(_06334_ ), .ZN(_06377_ ) );
XNOR2_X1 _14069_ ( .A(_06377_ ), .B(\u_lsu.u_clint.mtime [44] ), .ZN(_06378_ ) );
NOR2_X1 _14070_ ( .A1(_06378_ ), .A2(_06373_ ), .ZN(_00575_ ) );
AND3_X1 _14071_ ( .A1(_06318_ ), .A2(_01672_ ), .A3(_06319_ ), .ZN(_06379_ ) );
OAI21_X1 _14072_ ( .A(_05622_ ), .B1(_06379_ ), .B2(\u_lsu.u_clint.mtime [61] ), .ZN(_06380_ ) );
AND4_X1 _14073_ ( .A1(\u_lsu.u_clint.mtime [61] ), .A2(_06318_ ), .A3(_01672_ ), .A4(_06319_ ), .ZN(_06381_ ) );
NOR2_X1 _14074_ ( .A1(_06380_ ), .A2(_06381_ ), .ZN(_00576_ ) );
INV_X1 _14075_ ( .A(_06303_ ), .ZN(_06382_ ) );
NOR2_X1 _14076_ ( .A1(_06382_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ), .ZN(_06383_ ) );
AND2_X1 _14077_ ( .A1(_06383_ ), .A2(\u_lsu.u_clint.mtime [43] ), .ZN(_06384_ ) );
OAI21_X1 _14078_ ( .A(_04476_ ), .B1(_06383_ ), .B2(\u_lsu.u_clint.mtime [43] ), .ZN(_06385_ ) );
NOR2_X1 _14079_ ( .A1(_06384_ ), .A2(_06385_ ), .ZN(_00577_ ) );
AND3_X1 _14080_ ( .A1(_06333_ ), .A2(_06302_ ), .A3(_06369_ ), .ZN(_06386_ ) );
XNOR2_X1 _14081_ ( .A(_06386_ ), .B(\u_lsu.u_clint.mtime [42] ), .ZN(_06387_ ) );
NOR2_X1 _14082_ ( .A1(_06387_ ), .A2(_06373_ ), .ZN(_00578_ ) );
INV_X1 _14083_ ( .A(_06298_ ), .ZN(_06388_ ) );
INV_X1 _14084_ ( .A(_06300_ ), .ZN(_06389_ ) );
NOR3_X1 _14085_ ( .A1(_06388_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ), .A3(_06389_ ), .ZN(_06390_ ) );
OAI21_X1 _14086_ ( .A(_04473_ ), .B1(_06390_ ), .B2(\u_lsu.u_clint.mtime [41] ), .ZN(_06391_ ) );
AOI21_X1 _14087_ ( .A(_06391_ ), .B1(\u_lsu.u_clint.mtime [41] ), .B2(_06390_ ), .ZN(_00579_ ) );
XNOR2_X1 _14088_ ( .A(_06370_ ), .B(\u_lsu.u_clint.mtime [40] ), .ZN(_06392_ ) );
NOR2_X1 _14089_ ( .A1(_06392_ ), .A2(_06373_ ), .ZN(_00580_ ) );
NAND3_X1 _14090_ ( .A1(_06296_ ), .A2(\u_lsu.u_clint.mtime [36] ), .A3(_06297_ ), .ZN(_06393_ ) );
INV_X1 _14091_ ( .A(\u_lsu.u_clint.mtime [37] ), .ZN(_06394_ ) );
NOR3_X1 _14092_ ( .A1(_06393_ ), .A2(_06394_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ), .ZN(_06395_ ) );
AND2_X1 _14093_ ( .A1(_06395_ ), .A2(\u_lsu.u_clint.mtime [39] ), .ZN(_06396_ ) );
OAI21_X1 _14094_ ( .A(_04476_ ), .B1(_06395_ ), .B2(\u_lsu.u_clint.mtime [39] ), .ZN(_06397_ ) );
NOR2_X1 _14095_ ( .A1(_06396_ ), .A2(_06397_ ), .ZN(_00581_ ) );
AND3_X1 _14096_ ( .A1(_06333_ ), .A2(_06299_ ), .A3(_06335_ ), .ZN(_06398_ ) );
XNOR2_X1 _14097_ ( .A(_06398_ ), .B(\u_lsu.u_clint.mtime [38] ), .ZN(_06399_ ) );
NOR2_X1 _14098_ ( .A1(_06399_ ), .A2(_06373_ ), .ZN(_00582_ ) );
NAND3_X1 _14099_ ( .A1(_06296_ ), .A2(_02522_ ), .A3(_06297_ ), .ZN(_06400_ ) );
AOI21_X1 _14100_ ( .A(_02455_ ), .B1(_06400_ ), .B2(_06394_ ), .ZN(_06401_ ) );
NAND4_X1 _14101_ ( .A1(_06296_ ), .A2(\u_lsu.u_clint.mtime [37] ), .A3(_02522_ ), .A4(_06297_ ), .ZN(_06402_ ) );
AND2_X1 _14102_ ( .A1(_06401_ ), .A2(_06402_ ), .ZN(_00583_ ) );
AND2_X1 _14103_ ( .A1(_06333_ ), .A2(_06335_ ), .ZN(_06403_ ) );
XNOR2_X1 _14104_ ( .A(_06403_ ), .B(\u_lsu.u_clint.mtime [36] ), .ZN(_06404_ ) );
NOR2_X1 _14105_ ( .A1(_06404_ ), .A2(_06373_ ), .ZN(_00584_ ) );
NAND3_X1 _14106_ ( .A1(_06294_ ), .A2(_02626_ ), .A3(_06295_ ), .ZN(_06405_ ) );
AOI21_X1 _14107_ ( .A(_00893_ ), .B1(_06405_ ), .B2(_02576_ ), .ZN(_06406_ ) );
NAND4_X1 _14108_ ( .A1(_06294_ ), .A2(\u_lsu.u_clint.mtime [35] ), .A3(_02626_ ), .A4(_06295_ ), .ZN(_06407_ ) );
AND2_X1 _14109_ ( .A1(_06406_ ), .A2(_06407_ ), .ZN(_00585_ ) );
AND3_X1 _14110_ ( .A1(_06328_ ), .A2(_06295_ ), .A3(_06332_ ), .ZN(_06408_ ) );
XNOR2_X1 _14111_ ( .A(_06408_ ), .B(\u_lsu.u_clint.mtime [34] ), .ZN(_06409_ ) );
NOR2_X1 _14112_ ( .A1(_06409_ ), .A2(_06373_ ), .ZN(_00586_ ) );
XNOR2_X1 _14113_ ( .A(_06341_ ), .B(\u_lsu.u_clint.mtime [60] ), .ZN(_06410_ ) );
NOR2_X1 _14114_ ( .A1(_06410_ ), .A2(_06373_ ), .ZN(_00587_ ) );
AND3_X1 _14115_ ( .A1(_06292_ ), .A2(_02801_ ), .A3(_06293_ ), .ZN(_06411_ ) );
OAI21_X1 _14116_ ( .A(_05622_ ), .B1(_06411_ ), .B2(\u_lsu.u_clint.mtime [33] ), .ZN(_06412_ ) );
AND4_X1 _14117_ ( .A1(\u_lsu.u_clint.mtime [33] ), .A2(_06292_ ), .A3(_02801_ ), .A4(_06293_ ), .ZN(_06413_ ) );
NOR2_X1 _14118_ ( .A1(_06412_ ), .A2(_06413_ ), .ZN(_00588_ ) );
OR3_X1 _14119_ ( .A1(_06359_ ), .A2(\u_lsu.u_clint.mtime [32] ), .A3(_06360_ ), .ZN(_06414_ ) );
OAI21_X1 _14120_ ( .A(\u_lsu.u_clint.mtime [32] ), .B1(_06359_ ), .B2(_06360_ ), .ZN(_06415_ ) );
AOI211_X1 _14121_ ( .A(_05717_ ), .B(_00880_ ), .C1(_06414_ ), .C2(_06415_ ), .ZN(_00589_ ) );
AND2_X1 _14122_ ( .A1(_06328_ ), .A2(_06330_ ), .ZN(_06416_ ) );
NAND3_X1 _14123_ ( .A1(_06416_ ), .A2(_06291_ ), .A3(_06331_ ), .ZN(_06417_ ) );
NOR2_X1 _14124_ ( .A1(_06417_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_31_A_$_ANDNOT__Y_B ), .ZN(_06418_ ) );
XNOR2_X1 _14125_ ( .A(_06418_ ), .B(\u_lsu.u_clint.mtime [31] ), .ZN(_06419_ ) );
NOR2_X1 _14126_ ( .A1(_06419_ ), .A2(_06373_ ), .ZN(_00590_ ) );
OR2_X1 _14127_ ( .A1(_06417_ ), .A2(\u_lsu.u_clint.mtime [30] ), .ZN(_06420_ ) );
NAND2_X1 _14128_ ( .A1(_06417_ ), .A2(\u_lsu.u_clint.mtime [30] ), .ZN(_06421_ ) );
AOI21_X1 _14129_ ( .A(_00894_ ), .B1(_06420_ ), .B2(_06421_ ), .ZN(_00591_ ) );
AND2_X1 _14130_ ( .A1(_06416_ ), .A2(_06331_ ), .ZN(_06422_ ) );
INV_X1 _14131_ ( .A(_06422_ ), .ZN(_06423_ ) );
OR3_X1 _14132_ ( .A1(_06423_ ), .A2(\u_lsu.u_clint.mtime [29] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ), .ZN(_06424_ ) );
OAI21_X1 _14133_ ( .A(\u_lsu.u_clint.mtime [29] ), .B1(_06423_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ), .ZN(_06425_ ) );
AOI21_X1 _14134_ ( .A(_00894_ ), .B1(_06424_ ), .B2(_06425_ ), .ZN(_00592_ ) );
XNOR2_X1 _14135_ ( .A(_06422_ ), .B(\u_lsu.u_clint.mtime [28] ), .ZN(_06426_ ) );
NOR2_X1 _14136_ ( .A1(_06426_ ), .A2(_06373_ ), .ZN(_00593_ ) );
INV_X1 _14137_ ( .A(_06288_ ), .ZN(_06427_ ) );
NOR2_X1 _14138_ ( .A1(_06427_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ), .ZN(_06428_ ) );
OAI21_X1 _14139_ ( .A(_05622_ ), .B1(_06428_ ), .B2(\u_lsu.u_clint.mtime [27] ), .ZN(_06429_ ) );
NOR3_X1 _14140_ ( .A1(_06427_ ), .A2(_01731_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ), .ZN(_06430_ ) );
NOR2_X1 _14141_ ( .A1(_06429_ ), .A2(_06430_ ), .ZN(_00594_ ) );
AND3_X1 _14142_ ( .A1(_06328_ ), .A2(_06287_ ), .A3(_06330_ ), .ZN(_06431_ ) );
XNOR2_X1 _14143_ ( .A(_06431_ ), .B(\u_lsu.u_clint.mtime [26] ), .ZN(_06432_ ) );
NOR2_X1 _14144_ ( .A1(_06432_ ), .A2(_04470_ ), .ZN(_00595_ ) );
INV_X1 _14145_ ( .A(_06416_ ), .ZN(_06433_ ) );
OR3_X1 _14146_ ( .A1(_06433_ ), .A2(\u_lsu.u_clint.mtime [25] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ), .ZN(_06434_ ) );
OAI21_X1 _14147_ ( .A(\u_lsu.u_clint.mtime [25] ), .B1(_06433_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ), .ZN(_06435_ ) );
AOI21_X1 _14148_ ( .A(_00894_ ), .B1(_06434_ ), .B2(_06435_ ), .ZN(_00596_ ) );
XNOR2_X1 _14149_ ( .A(_06416_ ), .B(\u_lsu.u_clint.mtime [24] ), .ZN(_06436_ ) );
NOR2_X1 _14150_ ( .A1(_04461_ ), .A2(_06436_ ), .ZN(_00597_ ) );
AND3_X1 _14151_ ( .A1(_06316_ ), .A2(_01793_ ), .A3(_06317_ ), .ZN(_06437_ ) );
OAI21_X1 _14152_ ( .A(_05622_ ), .B1(_06437_ ), .B2(\u_lsu.u_clint.mtime [59] ), .ZN(_06438_ ) );
AND4_X1 _14153_ ( .A1(\u_lsu.u_clint.mtime [59] ), .A2(_06316_ ), .A3(_01793_ ), .A4(_06317_ ), .ZN(_06439_ ) );
NOR2_X1 _14154_ ( .A1(_06438_ ), .A2(_06439_ ), .ZN(_00598_ ) );
NAND3_X1 _14155_ ( .A1(_06328_ ), .A2(_06283_ ), .A3(_06329_ ), .ZN(_06440_ ) );
NOR2_X1 _14156_ ( .A1(_06440_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_39_A_$_ANDNOT__Y_B ), .ZN(_06441_ ) );
XNOR2_X1 _14157_ ( .A(_06441_ ), .B(\u_lsu.u_clint.mtime [23] ), .ZN(_06442_ ) );
NOR2_X1 _14158_ ( .A1(_06442_ ), .A2(_04470_ ), .ZN(_00599_ ) );
OR2_X1 _14159_ ( .A1(_06440_ ), .A2(\u_lsu.u_clint.mtime [22] ), .ZN(_06443_ ) );
NAND2_X1 _14160_ ( .A1(_06440_ ), .A2(\u_lsu.u_clint.mtime [22] ), .ZN(_06444_ ) );
AOI211_X1 _14161_ ( .A(_05717_ ), .B(_00880_ ), .C1(_06443_ ), .C2(_06444_ ), .ZN(_00600_ ) );
AND2_X1 _14162_ ( .A1(_06328_ ), .A2(_06329_ ), .ZN(_06445_ ) );
INV_X1 _14163_ ( .A(_06445_ ), .ZN(_06446_ ) );
OR3_X1 _14164_ ( .A1(_06446_ ), .A2(\u_lsu.u_clint.mtime [21] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ), .ZN(_06447_ ) );
OAI21_X1 _14165_ ( .A(\u_lsu.u_clint.mtime [21] ), .B1(_06446_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ), .ZN(_06448_ ) );
AOI21_X1 _14166_ ( .A(_00894_ ), .B1(_06447_ ), .B2(_06448_ ), .ZN(_00601_ ) );
AND4_X1 _14167_ ( .A1(\u_lsu.u_clint.mtime [11] ), .A2(_06272_ ), .A3(\u_lsu.u_clint.mtime [9] ), .A4(\u_lsu.u_clint.mtime [8] ), .ZN(_06449_ ) );
AND3_X1 _14168_ ( .A1(_06449_ ), .A2(\u_lsu.u_clint.mtime [13] ), .A3(\u_lsu.u_clint.mtime [10] ), .ZN(_06450_ ) );
AND3_X1 _14169_ ( .A1(_06450_ ), .A2(\u_lsu.u_clint.mtime [15] ), .A3(\u_lsu.u_clint.mtime [12] ), .ZN(_06451_ ) );
AND3_X1 _14170_ ( .A1(_06451_ ), .A2(\u_lsu.u_clint.mtime [17] ), .A3(\u_lsu.u_clint.mtime [14] ), .ZN(_06452_ ) );
AND2_X1 _14171_ ( .A1(_06452_ ), .A2(\u_lsu.u_clint.mtime [16] ), .ZN(_06453_ ) );
NAND4_X1 _14172_ ( .A1(_06453_ ), .A2(\u_lsu.u_clint.mtime [19] ), .A3(\u_lsu.u_clint.mtime [20] ), .A4(\u_lsu.u_clint.mtime [18] ), .ZN(_06454_ ) );
AND2_X1 _14173_ ( .A1(_06454_ ), .A2(_04473_ ), .ZN(_06455_ ) );
AND3_X1 _14174_ ( .A1(_06452_ ), .A2(\u_lsu.u_clint.mtime [19] ), .A3(\u_lsu.u_clint.mtime [16] ), .ZN(_06456_ ) );
AND2_X1 _14175_ ( .A1(_06456_ ), .A2(\u_lsu.u_clint.mtime [18] ), .ZN(_06457_ ) );
OAI21_X1 _14176_ ( .A(_06455_ ), .B1(\u_lsu.u_clint.mtime [20] ), .B2(_06457_ ), .ZN(_06458_ ) );
INV_X1 _14177_ ( .A(_06458_ ), .ZN(_00602_ ) );
INV_X1 _14178_ ( .A(_06280_ ), .ZN(_06459_ ) );
NOR2_X1 _14179_ ( .A1(_06459_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ), .ZN(_06460_ ) );
OAI21_X1 _14180_ ( .A(_04474_ ), .B1(_06460_ ), .B2(\u_lsu.u_clint.mtime [19] ), .ZN(_06461_ ) );
NOR3_X1 _14181_ ( .A1(_06459_ ), .A2(_01726_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ), .ZN(_06462_ ) );
NOR2_X1 _14182_ ( .A1(_06461_ ), .A2(_06462_ ), .ZN(_00603_ ) );
AND2_X1 _14183_ ( .A1(_06451_ ), .A2(\u_lsu.u_clint.mtime [14] ), .ZN(_06463_ ) );
NAND4_X1 _14184_ ( .A1(_06463_ ), .A2(\u_lsu.u_clint.mtime [17] ), .A3(\u_lsu.u_clint.mtime [18] ), .A4(\u_lsu.u_clint.mtime [16] ), .ZN(_06464_ ) );
AND2_X1 _14185_ ( .A1(_06464_ ), .A2(_04473_ ), .ZN(_06465_ ) );
OAI21_X1 _14186_ ( .A(_06465_ ), .B1(\u_lsu.u_clint.mtime [18] ), .B2(_06453_ ), .ZN(_06466_ ) );
INV_X1 _14187_ ( .A(_06466_ ), .ZN(_00604_ ) );
NOR4_X1 _14188_ ( .A1(_06325_ ), .A2(\u_lsu.u_clint.mtime [17] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ), .A4(_06327_ ), .ZN(_06467_ ) );
NOR3_X1 _14189_ ( .A1(_06325_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ), .A3(_06327_ ), .ZN(_06468_ ) );
NOR2_X1 _14190_ ( .A1(_06468_ ), .A2(_01879_ ), .ZN(_06469_ ) );
OAI211_X1 _14191_ ( .A(_04454_ ), .B(_00866_ ), .C1(_06467_ ), .C2(_06469_ ), .ZN(_06470_ ) );
INV_X1 _14192_ ( .A(_06470_ ), .ZN(_00605_ ) );
OAI21_X1 _14193_ ( .A(\u_lsu.u_clint.mtime [16] ), .B1(_06325_ ), .B2(_06327_ ), .ZN(_06471_ ) );
OR4_X1 _14194_ ( .A1(\u_lsu.u_clint.mtime [16] ), .A2(_06270_ ), .A3(_06327_ ), .A4(_06271_ ), .ZN(_06472_ ) );
AOI211_X1 _14195_ ( .A(_05717_ ), .B(_00880_ ), .C1(_06471_ ), .C2(_06472_ ), .ZN(_00606_ ) );
INV_X1 _14196_ ( .A(_06450_ ), .ZN(_06473_ ) );
INV_X1 _14197_ ( .A(\u_lsu.u_clint.mtime [12] ), .ZN(_06474_ ) );
NOR3_X1 _14198_ ( .A1(_06473_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ), .A3(_06474_ ), .ZN(_06475_ ) );
OAI21_X1 _14199_ ( .A(_04474_ ), .B1(_06475_ ), .B2(\u_lsu.u_clint.mtime [15] ), .ZN(_06476_ ) );
INV_X1 _14200_ ( .A(_06276_ ), .ZN(_06477_ ) );
NOR3_X1 _14201_ ( .A1(_06477_ ), .A2(_01231_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ), .ZN(_06478_ ) );
NOR2_X1 _14202_ ( .A1(_06476_ ), .A2(_06478_ ), .ZN(_00607_ ) );
AND2_X1 _14203_ ( .A1(_06449_ ), .A2(\u_lsu.u_clint.mtime [10] ), .ZN(_06479_ ) );
NAND4_X1 _14204_ ( .A1(_06479_ ), .A2(\u_lsu.u_clint.mtime [13] ), .A3(\u_lsu.u_clint.mtime [14] ), .A4(\u_lsu.u_clint.mtime [12] ), .ZN(_06480_ ) );
AND2_X1 _14205_ ( .A1(_04473_ ), .A2(_06480_ ), .ZN(_06481_ ) );
AND2_X1 _14206_ ( .A1(_06450_ ), .A2(\u_lsu.u_clint.mtime [12] ), .ZN(_06482_ ) );
OAI21_X1 _14207_ ( .A(_06481_ ), .B1(\u_lsu.u_clint.mtime [14] ), .B2(_06482_ ), .ZN(_06483_ ) );
INV_X1 _14208_ ( .A(_06483_ ), .ZN(_00608_ ) );
NAND3_X1 _14209_ ( .A1(_06337_ ), .A2(_06317_ ), .A3(_06338_ ), .ZN(_06484_ ) );
OR2_X1 _14210_ ( .A1(_06484_ ), .A2(\u_lsu.u_clint.mtime [58] ), .ZN(_06485_ ) );
NAND2_X1 _14211_ ( .A1(_06484_ ), .A2(\u_lsu.u_clint.mtime [58] ), .ZN(_06486_ ) );
AOI21_X1 _14212_ ( .A(_00894_ ), .B1(_06485_ ), .B2(_06486_ ), .ZN(_00609_ ) );
INV_X1 _14213_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ), .ZN(_06487_ ) );
AND3_X1 _14214_ ( .A1(_06274_ ), .A2(\u_lsu.u_clint.mtime [11] ), .A3(_06487_ ), .ZN(_06488_ ) );
OAI211_X1 _14215_ ( .A(_00863_ ), .B(_06068_ ), .C1(\u_lsu.u_clint.mtime [13] ), .C2(_06488_ ), .ZN(_06489_ ) );
AND4_X1 _14216_ ( .A1(\u_lsu.u_clint.mtime [13] ), .A2(_06274_ ), .A3(\u_lsu.u_clint.mtime [11] ), .A4(_06487_ ), .ZN(_06490_ ) );
OR2_X1 _14217_ ( .A1(_06489_ ), .A2(_06490_ ), .ZN(_06491_ ) );
INV_X1 _14218_ ( .A(_06491_ ), .ZN(_00610_ ) );
NAND3_X1 _14219_ ( .A1(_06449_ ), .A2(\u_lsu.u_clint.mtime [12] ), .A3(\u_lsu.u_clint.mtime [10] ), .ZN(_06492_ ) );
NAND3_X1 _14220_ ( .A1(_00863_ ), .A2(_06068_ ), .A3(_06492_ ), .ZN(_06493_ ) );
INV_X1 _14221_ ( .A(_06479_ ), .ZN(_06494_ ) );
AOI21_X1 _14222_ ( .A(_06493_ ), .B1(_06474_ ), .B2(_06494_ ), .ZN(_00611_ ) );
AND2_X1 _14223_ ( .A1(_06272_ ), .A2(_06273_ ), .ZN(_06495_ ) );
INV_X1 _14224_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ), .ZN(_06496_ ) );
AOI21_X1 _14225_ ( .A(\u_lsu.u_clint.mtime [11] ), .B1(_06495_ ), .B2(_06496_ ), .ZN(_06497_ ) );
AND4_X1 _14226_ ( .A1(\u_lsu.u_clint.mtime [11] ), .A2(_06272_ ), .A3(_06496_ ), .A4(_06273_ ), .ZN(_06498_ ) );
NOR4_X1 _14227_ ( .A1(flush_$_OR__Y_B ), .A2(_06497_ ), .A3(_05717_ ), .A4(_06498_ ), .ZN(_00612_ ) );
AOI21_X1 _14228_ ( .A(\u_lsu.u_clint.mtime [10] ), .B1(_06272_ ), .B2(_06273_ ), .ZN(_06499_ ) );
NOR4_X1 _14229_ ( .A1(flush_$_OR__Y_B ), .A2(_00882_ ), .A3(_06274_ ), .A4(_06499_ ), .ZN(_00613_ ) );
OR4_X1 _14230_ ( .A1(\u_lsu.u_clint.mtime [9] ), .A2(_06270_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ), .A4(_06271_ ), .ZN(_06500_ ) );
OAI21_X1 _14231_ ( .A(\u_lsu.u_clint.mtime [9] ), .B1(_06325_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ), .ZN(_06501_ ) );
AOI211_X1 _14232_ ( .A(_05717_ ), .B(_00880_ ), .C1(_06500_ ), .C2(_06501_ ), .ZN(_00614_ ) );
XNOR2_X1 _14233_ ( .A(_06272_ ), .B(\u_lsu.u_clint.mtime [8] ), .ZN(_06502_ ) );
NOR4_X1 _14234_ ( .A1(_04456_ ), .A2(_06502_ ), .A3(_06067_ ), .A4(reset ), .ZN(_00615_ ) );
OR3_X1 _14235_ ( .A1(_06270_ ), .A2(\u_lsu.u_clint.mtime [7] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ), .ZN(_06503_ ) );
OAI21_X1 _14236_ ( .A(\u_lsu.u_clint.mtime [7] ), .B1(_06270_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ), .ZN(_06504_ ) );
AOI211_X1 _14237_ ( .A(_05717_ ), .B(_00880_ ), .C1(_06503_ ), .C2(_06504_ ), .ZN(_00616_ ) );
XNOR2_X1 _14238_ ( .A(_06269_ ), .B(\u_lsu.u_clint.mtime [6] ), .ZN(_06505_ ) );
NOR4_X1 _14239_ ( .A1(_04456_ ), .A2(reset ), .A3(_06067_ ), .A4(_06505_ ), .ZN(_00617_ ) );
NOR3_X1 _14240_ ( .A1(_06266_ ), .A2(_02577_ ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ), .ZN(_06506_ ) );
XNOR2_X1 _14241_ ( .A(_06506_ ), .B(\u_lsu.u_clint.mtime [5] ), .ZN(_06507_ ) );
NOR4_X1 _14242_ ( .A1(_04456_ ), .A2(reset ), .A3(_06067_ ), .A4(_06507_ ), .ZN(_00618_ ) );
XNOR2_X1 _14243_ ( .A(_06267_ ), .B(\u_lsu.u_clint.mtime [4] ), .ZN(_06508_ ) );
NOR4_X1 _14244_ ( .A1(_04456_ ), .A2(reset ), .A3(_06067_ ), .A4(_06508_ ), .ZN(_00619_ ) );
INV_X1 _14245_ ( .A(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ), .ZN(_06509_ ) );
AND3_X1 _14246_ ( .A1(_06314_ ), .A2(_06509_ ), .A3(_06315_ ), .ZN(_06510_ ) );
OAI21_X1 _14247_ ( .A(_04474_ ), .B1(_06510_ ), .B2(\u_lsu.u_clint.mtime [57] ), .ZN(_06511_ ) );
AND4_X1 _14248_ ( .A1(\u_lsu.u_clint.mtime [57] ), .A2(_06314_ ), .A3(_06509_ ), .A4(_06315_ ), .ZN(_06512_ ) );
NOR2_X1 _14249_ ( .A1(_06511_ ), .A2(_06512_ ), .ZN(_00620_ ) );
AND2_X1 _14250_ ( .A1(\u_lsu.u_clint.mtime [1] ), .A2(\u_lsu.u_clint.mtime [0] ), .ZN(_06513_ ) );
INV_X1 _14251_ ( .A(_06513_ ), .ZN(_06514_ ) );
OR3_X1 _14252_ ( .A1(_06514_ ), .A2(\u_lsu.u_clint.mtime [3] ), .A3(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ), .ZN(_06515_ ) );
OAI21_X1 _14253_ ( .A(\u_lsu.u_clint.mtime [3] ), .B1(_06514_ ), .B2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ), .ZN(_06516_ ) );
AOI211_X1 _14254_ ( .A(_05717_ ), .B(_00880_ ), .C1(_06515_ ), .C2(_06516_ ), .ZN(_00621_ ) );
OR2_X1 _14255_ ( .A1(_06513_ ), .A2(\u_lsu.u_clint.mtime [2] ), .ZN(_06517_ ) );
AND4_X1 _14256_ ( .A1(_06061_ ), .A2(_00863_ ), .A3(_06266_ ), .A4(_06517_ ), .ZN(_00622_ ) );
NOR2_X1 _14257_ ( .A1(\u_lsu.u_clint.mtime [1] ), .A2(\u_lsu.u_clint.mtime [0] ), .ZN(_06518_ ) );
NOR4_X1 _14258_ ( .A1(_04455_ ), .A2(_00882_ ), .A3(_06513_ ), .A4(_06518_ ), .ZN(_00623_ ) );
AND3_X1 _14259_ ( .A1(_04454_ ), .A2(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D [0] ), .A3(_06061_ ), .ZN(_00624_ ) );
XNOR2_X1 _14260_ ( .A(_06339_ ), .B(\u_lsu.u_clint.mtime [56] ), .ZN(_06519_ ) );
NOR2_X1 _14261_ ( .A1(_06519_ ), .A2(_04470_ ), .ZN(_00625_ ) );
AND3_X1 _14262_ ( .A1(_06312_ ), .A2(_02000_ ), .A3(_06313_ ), .ZN(_06520_ ) );
OAI21_X1 _14263_ ( .A(_04474_ ), .B1(_06520_ ), .B2(\u_lsu.u_clint.mtime [55] ), .ZN(_06521_ ) );
AND4_X1 _14264_ ( .A1(\u_lsu.u_clint.mtime [55] ), .A2(_06312_ ), .A3(_02000_ ), .A4(_06313_ ), .ZN(_06522_ ) );
NOR2_X1 _14265_ ( .A1(_06521_ ), .A2(_06522_ ), .ZN(_00626_ ) );
NAND3_X1 _14266_ ( .A1(_06337_ ), .A2(_06313_ ), .A3(_06347_ ), .ZN(_06523_ ) );
OR2_X1 _14267_ ( .A1(_06523_ ), .A2(\u_lsu.u_clint.mtime [54] ), .ZN(_06524_ ) );
NAND2_X1 _14268_ ( .A1(_06523_ ), .A2(\u_lsu.u_clint.mtime [54] ), .ZN(_06525_ ) );
AOI21_X1 _14269_ ( .A(_00894_ ), .B1(_06524_ ), .B2(_06525_ ), .ZN(_00627_ ) );
INV_X1 _14270_ ( .A(\u_lsu.arvalid ), .ZN(_06526_ ) );
NOR4_X1 _14271_ ( .A1(_04456_ ), .A2(reset ), .A3(_06067_ ), .A4(_06526_ ), .ZN(_00628_ ) );
AND3_X1 _14272_ ( .A1(_00760_ ), .A2(\ea_errtp [0] ), .A3(ea_err ), .ZN(_00109_ ) );
NAND2_X1 _14273_ ( .A1(_01152_ ), .A2(_01154_ ), .ZN(\io_master_araddr [16] ) );
NAND2_X1 _14274_ ( .A1(_01153_ ), .A2(_01155_ ), .ZN(\io_master_araddr [23] ) );
NAND2_X1 _14275_ ( .A1(_01221_ ), .A2(_01222_ ), .ZN(\io_master_araddr [8] ) );
NOR2_X1 _14276_ ( .A1(_01173_ ), .A2(_01172_ ), .ZN(\io_master_araddr [14] ) );
INV_X1 _14277_ ( .A(_01239_ ), .ZN(\io_master_araddr [2] ) );
AND2_X1 _14278_ ( .A1(_01275_ ), .A2(\u_arbiter.rmask [1] ), .ZN(\io_master_arsize [0] ) );
NOR2_X1 _14279_ ( .A1(_01909_ ), .A2(_06526_ ), .ZN(io_master_arvalid ) );
NAND2_X1 _14280_ ( .A1(io_master_awready ), .A2(io_master_awvalid ), .ZN(_06527_ ) );
OAI21_X1 _14281_ ( .A(_06527_ ), .B1(_06249_ ), .B2(\u_lsu.writing ), .ZN(\u_lsu.awvalid_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14282_ ( .A(\al_wmask [1] ), .ZN(_06528_ ) );
NOR2_X1 _14283_ ( .A1(_06528_ ), .A2(\al_wmask [0] ), .ZN(\io_master_awsize [0] ) );
AND2_X1 _14284_ ( .A1(\al_wmask [1] ), .A2(\al_wmask [0] ), .ZN(\io_master_awsize [1] ) );
NOR2_X1 _14285_ ( .A1(_06249_ ), .A2(\u_lsu.writing ), .ZN(_06529_ ) );
OR2_X1 _14286_ ( .A1(_06529_ ), .A2(io_master_bvalid ), .ZN(io_master_bvalid_$_OR__B_Y ) );
INV_X1 _14287_ ( .A(\al_wdata [7] ), .ZN(_06530_ ) );
NOR3_X1 _14288_ ( .A1(_06530_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [7] ) );
INV_X1 _14289_ ( .A(\al_wdata [6] ), .ZN(_06531_ ) );
NOR3_X1 _14290_ ( .A1(_06531_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [6] ) );
INV_X1 _14291_ ( .A(\al_wdata [5] ), .ZN(_06532_ ) );
NOR3_X1 _14292_ ( .A1(_06532_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [5] ) );
INV_X1 _14293_ ( .A(\al_wdata [4] ), .ZN(_06533_ ) );
NOR3_X1 _14294_ ( .A1(_06533_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [4] ) );
INV_X1 _14295_ ( .A(\al_wdata [3] ), .ZN(_06534_ ) );
NOR3_X1 _14296_ ( .A1(_06534_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14297_ ( .A(\al_wdata [2] ), .ZN(_06535_ ) );
NOR3_X1 _14298_ ( .A1(_06535_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14299_ ( .A(\al_wdata [1] ), .ZN(_06536_ ) );
NOR3_X1 _14300_ ( .A1(_06536_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14301_ ( .A(\al_wdata [0] ), .ZN(_06537_ ) );
NOR3_X1 _14302_ ( .A1(_06537_ ), .A2(\io_master_awaddr [0] ), .A3(\io_master_awaddr [1] ), .ZN(\io_master_wdata [0] ) );
INV_X1 _14303_ ( .A(\io_master_awaddr [0] ), .ZN(_06538_ ) );
NOR2_X1 _14304_ ( .A1(_06538_ ), .A2(\io_master_awaddr [1] ), .ZN(_06539_ ) );
NOR2_X1 _14305_ ( .A1(\io_master_awaddr [0] ), .A2(\io_master_awaddr [1] ), .ZN(_06540_ ) );
AOI22_X1 _14306_ ( .A1(_06539_ ), .A2(\al_wdata [23] ), .B1(_06540_ ), .B2(\al_wdata [31] ), .ZN(_06541_ ) );
AND2_X1 _14307_ ( .A1(\io_master_awaddr [0] ), .A2(\io_master_awaddr [1] ), .ZN(_06542_ ) );
INV_X1 _14308_ ( .A(_06542_ ), .ZN(_06543_ ) );
INV_X1 _14309_ ( .A(\al_wdata [15] ), .ZN(_06544_ ) );
INV_X1 _14310_ ( .A(\io_master_awaddr [1] ), .ZN(_06545_ ) );
NOR2_X1 _14311_ ( .A1(_06545_ ), .A2(\io_master_awaddr [0] ), .ZN(_06546_ ) );
INV_X1 _14312_ ( .A(_06546_ ), .ZN(_06547_ ) );
BUF_X4 _14313_ ( .A(_06547_ ), .Z(_06548_ ) );
OAI221_X1 _14314_ ( .A(_06541_ ), .B1(_06530_ ), .B2(_06543_ ), .C1(_06544_ ), .C2(_06548_ ), .ZN(\io_master_wdata [31] ) );
AOI22_X1 _14315_ ( .A1(_06546_ ), .A2(\al_wdata [14] ), .B1(_06540_ ), .B2(\al_wdata [30] ), .ZN(_06549_ ) );
INV_X1 _14316_ ( .A(\al_wdata [22] ), .ZN(_06550_ ) );
INV_X2 _14317_ ( .A(_06539_ ), .ZN(_06551_ ) );
OAI221_X1 _14318_ ( .A(_06549_ ), .B1(_06531_ ), .B2(_06543_ ), .C1(_06550_ ), .C2(_06551_ ), .ZN(\io_master_wdata [30] ) );
BUF_X4 _14319_ ( .A(_06538_ ), .Z(_06552_ ) );
BUF_X4 _14320_ ( .A(_06545_ ), .Z(_06553_ ) );
NAND3_X1 _14321_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [21] ), .ZN(_06554_ ) );
INV_X1 _14322_ ( .A(\al_wdata [13] ), .ZN(_06555_ ) );
OAI221_X1 _14323_ ( .A(_06554_ ), .B1(_06548_ ), .B2(_06532_ ), .C1(_06555_ ), .C2(_06551_ ), .ZN(\io_master_wdata [21] ) );
NAND3_X1 _14324_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [20] ), .ZN(_06556_ ) );
INV_X1 _14325_ ( .A(\al_wdata [12] ), .ZN(_06557_ ) );
OAI221_X1 _14326_ ( .A(_06556_ ), .B1(_06548_ ), .B2(_06533_ ), .C1(_06557_ ), .C2(_06551_ ), .ZN(\io_master_wdata [20] ) );
NAND3_X1 _14327_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [19] ), .ZN(_06558_ ) );
INV_X1 _14328_ ( .A(\al_wdata [11] ), .ZN(_06559_ ) );
OAI221_X1 _14329_ ( .A(_06558_ ), .B1(_06548_ ), .B2(_06534_ ), .C1(_06559_ ), .C2(_06551_ ), .ZN(\io_master_wdata [19] ) );
NAND3_X1 _14330_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [18] ), .ZN(_06560_ ) );
INV_X1 _14331_ ( .A(\al_wdata [10] ), .ZN(_06561_ ) );
OAI221_X1 _14332_ ( .A(_06560_ ), .B1(_06548_ ), .B2(_06535_ ), .C1(_06561_ ), .C2(_06551_ ), .ZN(\io_master_wdata [18] ) );
NAND3_X1 _14333_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [17] ), .ZN(_06562_ ) );
INV_X1 _14334_ ( .A(\al_wdata [9] ), .ZN(_06563_ ) );
OAI221_X1 _14335_ ( .A(_06562_ ), .B1(_06547_ ), .B2(_06536_ ), .C1(_06563_ ), .C2(_06551_ ), .ZN(\io_master_wdata [17] ) );
NAND3_X1 _14336_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [16] ), .ZN(_06564_ ) );
INV_X1 _14337_ ( .A(\al_wdata [8] ), .ZN(_06565_ ) );
OAI221_X1 _14338_ ( .A(_06564_ ), .B1(_06547_ ), .B2(_06537_ ), .C1(_06565_ ), .C2(_06551_ ), .ZN(\io_master_wdata [16] ) );
BUF_X4 _14339_ ( .A(_06551_ ), .Z(_06566_ ) );
INV_X2 _14340_ ( .A(_06540_ ), .ZN(_06567_ ) );
OAI22_X1 _14341_ ( .A1(_06566_ ), .A2(_06530_ ), .B1(_06544_ ), .B2(_06567_ ), .ZN(\io_master_wdata [15] ) );
INV_X1 _14342_ ( .A(\al_wdata [14] ), .ZN(_06568_ ) );
OAI22_X1 _14343_ ( .A1(_06566_ ), .A2(_06531_ ), .B1(_06568_ ), .B2(_06567_ ), .ZN(\io_master_wdata [14] ) );
OAI22_X1 _14344_ ( .A1(_06566_ ), .A2(_06532_ ), .B1(_06555_ ), .B2(_06567_ ), .ZN(\io_master_wdata [13] ) );
OAI22_X1 _14345_ ( .A1(_06566_ ), .A2(_06533_ ), .B1(_06557_ ), .B2(_06567_ ), .ZN(\io_master_wdata [12] ) );
AOI22_X1 _14346_ ( .A1(_06539_ ), .A2(\al_wdata [21] ), .B1(_06540_ ), .B2(\al_wdata [29] ), .ZN(_06569_ ) );
OAI221_X1 _14347_ ( .A(_06569_ ), .B1(_06532_ ), .B2(_06543_ ), .C1(_06555_ ), .C2(_06548_ ), .ZN(\io_master_wdata [29] ) );
OAI22_X1 _14348_ ( .A1(_06566_ ), .A2(_06534_ ), .B1(_06559_ ), .B2(_06567_ ), .ZN(\io_master_wdata [11] ) );
OAI22_X1 _14349_ ( .A1(_06566_ ), .A2(_06535_ ), .B1(_06561_ ), .B2(_06567_ ), .ZN(\io_master_wdata [10] ) );
OAI22_X1 _14350_ ( .A1(_06566_ ), .A2(_06536_ ), .B1(_06563_ ), .B2(_06567_ ), .ZN(\io_master_wdata [9] ) );
OAI22_X1 _14351_ ( .A1(_06566_ ), .A2(_06537_ ), .B1(_06565_ ), .B2(_06567_ ), .ZN(\io_master_wdata [8] ) );
AOI22_X1 _14352_ ( .A1(_06539_ ), .A2(\al_wdata [20] ), .B1(_06542_ ), .B2(\al_wdata [4] ), .ZN(_06570_ ) );
NAND3_X1 _14353_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [28] ), .ZN(_06571_ ) );
OAI211_X1 _14354_ ( .A(_06570_ ), .B(_06571_ ), .C1(_06557_ ), .C2(_06548_ ), .ZN(\io_master_wdata [28] ) );
AOI22_X1 _14355_ ( .A1(_06539_ ), .A2(\al_wdata [19] ), .B1(_06540_ ), .B2(\al_wdata [27] ), .ZN(_06572_ ) );
OAI221_X1 _14356_ ( .A(_06572_ ), .B1(_06534_ ), .B2(_06543_ ), .C1(_06559_ ), .C2(_06548_ ), .ZN(\io_master_wdata [27] ) );
AOI22_X1 _14357_ ( .A1(_06539_ ), .A2(\al_wdata [18] ), .B1(_06540_ ), .B2(\al_wdata [26] ), .ZN(_06573_ ) );
OAI221_X1 _14358_ ( .A(_06573_ ), .B1(_06535_ ), .B2(_06543_ ), .C1(_06561_ ), .C2(_06548_ ), .ZN(\io_master_wdata [26] ) );
AOI22_X1 _14359_ ( .A1(\al_wdata [17] ), .A2(_06539_ ), .B1(_06546_ ), .B2(\al_wdata [9] ), .ZN(_06574_ ) );
NAND3_X1 _14360_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [25] ), .ZN(_06575_ ) );
OAI211_X1 _14361_ ( .A(_06574_ ), .B(_06575_ ), .C1(_06536_ ), .C2(_06543_ ), .ZN(\io_master_wdata [25] ) );
AOI22_X1 _14362_ ( .A1(\al_wdata [16] ), .A2(_06539_ ), .B1(_06546_ ), .B2(\al_wdata [8] ), .ZN(_06576_ ) );
NAND3_X1 _14363_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [24] ), .ZN(_06577_ ) );
OAI211_X1 _14364_ ( .A(_06576_ ), .B(_06577_ ), .C1(_06537_ ), .C2(_06543_ ), .ZN(\io_master_wdata [24] ) );
NAND3_X1 _14365_ ( .A1(_06552_ ), .A2(_06553_ ), .A3(\al_wdata [23] ), .ZN(_06578_ ) );
OAI221_X1 _14366_ ( .A(_06578_ ), .B1(_06547_ ), .B2(_06530_ ), .C1(_06544_ ), .C2(_06551_ ), .ZN(\io_master_wdata [23] ) );
NAND3_X1 _14367_ ( .A1(_06538_ ), .A2(\al_wdata [6] ), .A3(\io_master_awaddr [1] ), .ZN(_06579_ ) );
OAI221_X1 _14368_ ( .A(_06579_ ), .B1(_06567_ ), .B2(_06550_ ), .C1(_06566_ ), .C2(_06568_ ), .ZN(\io_master_wdata [22] ) );
NAND2_X1 _14369_ ( .A1(io_master_wready ), .A2(io_master_wlast ), .ZN(_06580_ ) );
OAI21_X1 _14370_ ( .A(_06580_ ), .B1(_06249_ ), .B2(\u_lsu.writing ), .ZN(\u_lsu.wlast_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14371_ ( .A(\al_wmask [0] ), .ZN(_06581_ ) );
AND3_X1 _14372_ ( .A1(_06581_ ), .A2(\al_wmask [1] ), .A3(\io_master_awaddr [1] ), .ZN(_06582_ ) );
NOR2_X1 _14373_ ( .A1(_06582_ ), .A2(\io_master_awsize [1] ), .ZN(_06583_ ) );
OAI21_X1 _14374_ ( .A(_06583_ ), .B1(_06581_ ), .B2(_06543_ ), .ZN(\io_master_wstrb [3] ) );
OAI21_X1 _14375_ ( .A(_06583_ ), .B1(_06581_ ), .B2(_06548_ ), .ZN(\io_master_wstrb [2] ) );
NOR3_X1 _14376_ ( .A1(_06528_ ), .A2(\al_wmask [0] ), .A3(\io_master_awaddr [1] ), .ZN(_06584_ ) );
NOR2_X1 _14377_ ( .A1(_06584_ ), .A2(\io_master_awsize [1] ), .ZN(_06585_ ) );
OAI21_X1 _14378_ ( .A(_06585_ ), .B1(_06581_ ), .B2(_06566_ ), .ZN(\io_master_wstrb [1] ) );
OAI21_X1 _14379_ ( .A(_06585_ ), .B1(_06581_ ), .B2(_06567_ ), .ZN(\io_master_wstrb [0] ) );
NAND2_X1 _14380_ ( .A1(_00760_ ), .A2(_00777_ ), .ZN(_06586_ ) );
OAI22_X1 _14381_ ( .A1(_06047_ ), .A2(_01280_ ), .B1(_00762_ ), .B2(_06586_ ), .ZN(\u_arbiter.rvalid_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14382_ ( .A1(\u_lsu.writing ), .A2(io_master_bvalid ), .ZN(_06587_ ) );
OR2_X1 _14383_ ( .A1(_06249_ ), .A2(_06587_ ), .ZN(_06588_ ) );
NAND4_X1 _14384_ ( .A1(_01283_ ), .A2(_06586_ ), .A3(_01284_ ), .A4(_06588_ ), .ZN(\u_arbiter.working_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14385_ ( .A(_06588_ ), .B1(_06586_ ), .B2(\u_exu.eopt [12] ), .ZN(\u_arbiter.wvalid_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _14386_ ( .A1(_01384_ ), .A2(_01388_ ), .A3(_01430_ ), .ZN(_06589_ ) );
NAND2_X1 _14387_ ( .A1(_06589_ ), .A2(_01434_ ), .ZN(_06590_ ) );
NOR3_X1 _14388_ ( .A1(_06590_ ), .A2(_01391_ ), .A3(_01396_ ), .ZN(_06591_ ) );
NOR2_X1 _14389_ ( .A1(_01413_ ), .A2(_01399_ ), .ZN(_06592_ ) );
AND3_X1 _14390_ ( .A1(_06592_ ), .A2(_01411_ ), .A3(_01405_ ), .ZN(_06593_ ) );
AND4_X1 _14391_ ( .A1(_01427_ ), .A2(_06591_ ), .A3(_01377_ ), .A4(_06593_ ), .ZN(_06594_ ) );
AND2_X1 _14392_ ( .A1(_06594_ ), .A2(_01381_ ), .ZN(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _14393_ ( .A1(_01376_ ), .A2(_01427_ ), .ZN(_06595_ ) );
NAND3_X1 _14394_ ( .A1(_06595_ ), .A2(_01390_ ), .A3(_01396_ ), .ZN(_06596_ ) );
NOR2_X1 _14395_ ( .A1(_06590_ ), .A2(_06596_ ), .ZN(_06597_ ) );
AND4_X1 _14396_ ( .A1(_00760_ ), .A2(_06597_ ), .A3(_01380_ ), .A4(_06593_ ), .ZN(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y ) );
AND3_X1 _14397_ ( .A1(_06592_ ), .A2(_01411_ ), .A3(_01406_ ), .ZN(_06598_ ) );
AND4_X1 _14398_ ( .A1(_01381_ ), .A2(_06591_ ), .A3(_06595_ ), .A4(_06598_ ), .ZN(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OAI21_X1 _14399_ ( .A(_04485_ ), .B1(_00633_ ), .B2(_00636_ ), .ZN(\u_exu.exe_end_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14400_ ( .A(_01057_ ), .B1(_04484_ ), .B2(_00761_ ), .ZN(\u_exu.exe_start_$_SDFFE_PP0P__Q_E ) );
OR2_X1 _14401_ ( .A1(icah_ready ), .A2(_05547_ ), .ZN(\u_icache.caddr_$_SDFFE_PP0P__Q_E ) );
BUF_X4 _14402_ ( .A(_06048_ ), .Z(_06599_ ) );
NOR2_X1 _14403_ ( .A1(_01279_ ), .A2(_06599_ ), .ZN(\ac_data [31] ) );
NOR2_X1 _14404_ ( .A1(_01533_ ), .A2(_06599_ ), .ZN(\ac_data [30] ) );
NOR2_X1 _14405_ ( .A1(_01618_ ), .A2(_06599_ ), .ZN(\ac_data [21] ) );
NOR2_X1 _14406_ ( .A1(_01685_ ), .A2(_06599_ ), .ZN(\ac_data [20] ) );
NOR2_X1 _14407_ ( .A1(_01740_ ), .A2(_06599_ ), .ZN(\ac_data [19] ) );
NOR2_X1 _14408_ ( .A1(_01803_ ), .A2(_06599_ ), .ZN(\ac_data [18] ) );
NOR2_X1 _14409_ ( .A1(_01889_ ), .A2(_06599_ ), .ZN(\ac_data [17] ) );
NOR2_X1 _14410_ ( .A1(_01921_ ), .A2(_06599_ ), .ZN(\ac_data [16] ) );
NOR2_X1 _14411_ ( .A1(_01959_ ), .A2(_06599_ ), .ZN(\ac_data [15] ) );
NOR2_X1 _14412_ ( .A1(_02010_ ), .A2(_06599_ ), .ZN(\ac_data [14] ) );
BUF_X4 _14413_ ( .A(_06048_ ), .Z(_06600_ ) );
NOR2_X1 _14414_ ( .A1(_02063_ ), .A2(_06600_ ), .ZN(\ac_data [13] ) );
NOR2_X1 _14415_ ( .A1(_02107_ ), .A2(_06600_ ), .ZN(\ac_data [12] ) );
NOR2_X1 _14416_ ( .A1(_02145_ ), .A2(_06600_ ), .ZN(\ac_data [29] ) );
NOR2_X1 _14417_ ( .A1(_02189_ ), .A2(_06600_ ), .ZN(\ac_data [11] ) );
NOR2_X1 _14418_ ( .A1(_02235_ ), .A2(_06600_ ), .ZN(\ac_data [10] ) );
NOR2_X1 _14419_ ( .A1(_01604_ ), .A2(_02283_ ), .ZN(_06601_ ) );
NOR2_X1 _14420_ ( .A1(_06601_ ), .A2(_06600_ ), .ZN(\ac_data [9] ) );
NOR2_X1 _14421_ ( .A1(_02326_ ), .A2(_06600_ ), .ZN(\ac_data [8] ) );
OAI211_X1 _14422_ ( .A(_05551_ ), .B(_02431_ ), .C1(_01253_ ), .C2(_01258_ ), .ZN(_06602_ ) );
INV_X1 _14423_ ( .A(_06602_ ), .ZN(\ac_data [7] ) );
OAI211_X1 _14424_ ( .A(_05551_ ), .B(_02431_ ), .C1(_02434_ ), .C2(_02438_ ), .ZN(_06603_ ) );
INV_X1 _14425_ ( .A(_06603_ ), .ZN(\ac_data [6] ) );
AND4_X1 _14426_ ( .A1(_05551_ ), .A2(_02464_ ), .A3(_02431_ ), .A4(_02468_ ), .ZN(\ac_data [5] ) );
NAND2_X1 _14427_ ( .A1(_02527_ ), .A2(_05551_ ), .ZN(_06604_ ) );
INV_X1 _14428_ ( .A(_06604_ ), .ZN(\ac_data [4] ) );
AND4_X1 _14429_ ( .A1(_05551_ ), .A2(_02574_ ), .A3(_02431_ ), .A4(_02579_ ), .ZN(\ac_data [3] ) );
NAND2_X1 _14430_ ( .A1(_02631_ ), .A2(_05551_ ), .ZN(_06605_ ) );
INV_X1 _14431_ ( .A(_06605_ ), .ZN(\ac_data [2] ) );
NOR2_X1 _14432_ ( .A1(_02706_ ), .A2(_06600_ ), .ZN(\ac_data [28] ) );
AND4_X1 _14433_ ( .A1(_05551_ ), .A2(_02728_ ), .A3(_02431_ ), .A4(_02732_ ), .ZN(\ac_data [1] ) );
OAI211_X1 _14434_ ( .A(_05551_ ), .B(_02431_ ), .C1(_02804_ ), .C2(_02807_ ), .ZN(_06606_ ) );
INV_X1 _14435_ ( .A(_06606_ ), .ZN(\ac_data [0] ) );
NOR2_X1 _14436_ ( .A1(_02834_ ), .A2(_06600_ ), .ZN(\ac_data [27] ) );
NOR2_X1 _14437_ ( .A1(_02889_ ), .A2(_06600_ ), .ZN(\ac_data [26] ) );
NOR2_X1 _14438_ ( .A1(_02909_ ), .A2(_06048_ ), .ZN(\ac_data [25] ) );
NOR2_X1 _14439_ ( .A1(_02943_ ), .A2(_06048_ ), .ZN(\ac_data [24] ) );
NOR2_X1 _14440_ ( .A1(_03015_ ), .A2(_06048_ ), .ZN(\ac_data [23] ) );
NOR2_X1 _14441_ ( .A1(_03038_ ), .A2(_06048_ ), .ZN(\ac_data [22] ) );
NAND2_X1 _14442_ ( .A1(\fc_addr [4] ), .A2(\u_icache.count [1] ), .ZN(_06607_ ) );
NOR4_X1 _14443_ ( .A1(_06047_ ), .A2(\u_icache.count_$_NOT__A_Y ), .A3(_06048_ ), .A4(_06607_ ), .ZN(\u_icache.count_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14444_ ( .A1(_06045_ ), .A2(_05690_ ), .A3(\u_icache.count [1] ), .A4(\u_icache.count_$_NOT__A_Y ), .ZN(\u_icache.count_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _14445_ ( .A(\u_icache.count [1] ), .ZN(_06608_ ) );
NOR4_X1 _14446_ ( .A1(_06045_ ), .A2(\fc_addr [4] ), .A3(_06608_ ), .A4(\u_icache.count_$_NOT__A_Y ), .ZN(\u_icache.count_$_ORNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14447_ ( .A1(_06045_ ), .A2(\fc_addr [4] ), .A3(\u_icache.count [1] ), .A4(\u_icache.count_$_NOT__A_Y ), .ZN(\u_icache.count_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14448_ ( .A1(_06045_ ), .A2(\fc_addr [4] ), .A3(\u_icache.count [1] ), .A4(\u_icache.count [0] ), .ZN(\u_icache.count_$_OR__B_1_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14449_ ( .A1(_06045_ ), .A2(\fc_addr [4] ), .A3(_06608_ ), .A4(\u_icache.count [0] ), .ZN(\u_icache.count_$_OR__B_2_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14450_ ( .A1(_06047_ ), .A2(\u_icache.count [0] ), .A3(_06048_ ), .A4(_06607_ ), .ZN(\u_icache.count_$_OR__B_3_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14451_ ( .A1(_06045_ ), .A2(_05690_ ), .A3(\u_icache.count [1] ), .A4(\u_icache.count [0] ), .ZN(\u_icache.count_$_OR__B_Y_$_ANDNOT__B_Y ) );
OAI21_X1 _14452_ ( .A(_06052_ ), .B1(_06047_ ), .B2(_06048_ ), .ZN(\u_icache.count_$_SDFFE_PP0P__Q_E ) );
NAND3_X1 _14453_ ( .A1(icah_ready ), .A2(_06043_ ), .A3(_06042_ ), .ZN(_06609_ ) );
OAI21_X1 _14454_ ( .A(_06609_ ), .B1(_06049_ ), .B2(_05403_ ), .ZN(\u_icache.ended_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14455_ ( .A1(_06609_ ), .A2(_05698_ ), .ZN(\u_icache.chvalid_$_SDFFE_PP0P__Q_E ) );
OR2_X1 _14456_ ( .A1(_01090_ ), .A2(\u_exu.exe_end_$_ANDNOT__B_Y ), .ZN(\u_exu.alu_p2_$_SDFFE_PP0P__Q_E ) );
OR2_X1 _14457_ ( .A1(_01090_ ), .A2(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .ZN(\u_idu.decode_ok_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14458_ ( .A(_06055_ ), .B1(_05403_ ), .B2(_06049_ ), .ZN(\u_ifu.inst_ok_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _14459_ ( .A1(_05403_ ), .A2(_06049_ ), .B1(_00765_ ), .B2(_00759_ ), .ZN(\u_ifu.jpc_ok_$_SDFFE_PP0P__Q_E ) );
NOR4_X1 _14460_ ( .A1(_04456_ ), .A2(reset ), .A3(_06187_ ), .A4(_06052_ ), .ZN(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_Y ) );
NOR4_X1 _14461_ ( .A1(_04456_ ), .A2(reset ), .A3(_05690_ ), .A4(_06052_ ), .ZN(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_B_$_ANDNOT__B_Y ) );
MUX2_X1 _14462_ ( .A(_00858_ ), .B(_00766_ ), .S(_06130_ ), .Z(\u_ifu.pc_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14463_ ( .A(\u_lsu.arvalid ), .B1(_01909_ ), .B2(io_master_arready ), .ZN(_06610_ ) );
NAND2_X1 _14464_ ( .A1(_06610_ ), .A2(_06248_ ), .ZN(\u_lsu.arvalid_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14465_ ( .A1(\u_lsu.rvalid ), .A2(_06265_ ), .ZN(_06611_ ) );
NAND2_X1 _14466_ ( .A1(_06611_ ), .A2(_06248_ ), .ZN(\u_lsu.reading_$_SDFFE_PP0P__Q_E ) );
CLKGATE_X1 _14467_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_06612_ ) );
CLKGATE_X1 _14468_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_1_Y_$_ANDNOT__B_Y ), .GCK(_06613_ ) );
CLKGATE_X1 _14469_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_06614_ ) );
CLKGATE_X1 _14470_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06615_ ) );
CLKGATE_X1 _14471_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06616_ ) );
CLKGATE_X1 _14472_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ANDNOT__A_1_Y_$_AND__B_Y ), .GCK(_06617_ ) );
CLKGATE_X1 _14473_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .GCK(_06618_ ) );
CLKGATE_X1 _14474_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_06619_ ) );
CLKGATE_X1 _14475_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .GCK(_06620_ ) );
CLKGATE_X1 _14476_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06621_ ) );
CLKGATE_X1 _14477_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_1_Y_$_ANDNOT__B_Y ), .GCK(_06622_ ) );
CLKGATE_X1 _14478_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_6_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_06623_ ) );
CLKGATE_X1 _14479_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B_$_ORNOT__B_Y_$_ANDNOT__B_Y ), .GCK(_06624_ ) );
CLKGATE_X1 _14480_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_06625_ ) );
CLKGATE_X1 _14481_ ( .CK(clock ), .E(\u_exu.rlock_nxt_$_MUX__Y_5_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_06626_ ) );
CLKGATE_X1 _14482_ ( .CK(clock ), .E(io_master_bvalid_$_OR__B_Y ), .GCK(_06627_ ) );
CLKGATE_X1 _14483_ ( .CK(clock ), .E(\u_lsu.wlast_$_SDFFE_PP0P__Q_E ), .GCK(_06628_ ) );
CLKGATE_X1 _14484_ ( .CK(clock ), .E(\u_lsu.reading_$_SDFFE_PP0P__Q_E ), .GCK(_06629_ ) );
CLKGATE_X1 _14485_ ( .CK(clock ), .E(\u_lsu.rvalid ), .GCK(_06630_ ) );
CLKGATE_X1 _14486_ ( .CK(clock ), .E(\u_lsu.awvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06631_ ) );
CLKGATE_X1 _14487_ ( .CK(clock ), .E(\u_lsu.arvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06632_ ) );
CLKGATE_X1 _14488_ ( .CK(clock ), .E(\u_ifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_06633_ ) );
CLKGATE_X1 _14489_ ( .CK(clock ), .E(_00000_ ), .GCK(_06634_ ) );
CLKGATE_X1 _14490_ ( .CK(clock ), .E(\u_ifu.jpc_ok_$_SDFFE_PP0P__Q_E ), .GCK(_06635_ ) );
CLKGATE_X1 _14491_ ( .CK(clock ), .E(\u_ifu.inst_ok_$_SDFFE_PP0P__Q_E ), .GCK(_06636_ ) );
CLKGATE_X1 _14492_ ( .CK(clock ), .E(\u_icache.cready_$_ANDNOT__A_Y ), .GCK(_06637_ ) );
CLKGATE_X1 _14493_ ( .CK(clock ), .E(\u_ifu.inst_ok_$_ANDNOT__A_Y ), .GCK(_06638_ ) );
CLKGATE_X1 _14494_ ( .CK(clock ), .E(\u_idu.decode_ok_$_SDFFE_PP0P__Q_E ), .GCK(_06639_ ) );
CLKGATE_X1 _14495_ ( .CK(clock ), .E(\u_icache.ended_$_SDFFE_PP0P__Q_E ), .GCK(_06640_ ) );
CLKGATE_X1 _14496_ ( .CK(clock ), .E(\u_icache.cvalids_$_SDFFE_PP0P__Q_E ), .GCK(_06641_ ) );
CLKGATE_X1 _14497_ ( .CK(clock ), .E(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_B_$_ANDNOT__B_Y ), .GCK(_06642_ ) );
CLKGATE_X1 _14498_ ( .CK(clock ), .E(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__A_Y ), .GCK(_06643_ ) );
CLKGATE_X1 _14499_ ( .CK(clock ), .E(\u_icache.count_$_SDFFE_PP0P__Q_E ), .GCK(_06644_ ) );
CLKGATE_X1 _14500_ ( .CK(clock ), .E(\u_icache.chvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06645_ ) );
CLKGATE_X1 _14501_ ( .CK(clock ), .E(\u_icache.cready_$_ANDNOT__B_Y_$_OR__B_Y ), .GCK(_06646_ ) );
CLKGATE_X1 _14502_ ( .CK(clock ), .E(\u_icache.count_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06647_ ) );
CLKGATE_X1 _14503_ ( .CK(clock ), .E(\u_icache.count_$_OR__B_3_Y_$_ANDNOT__B_Y ), .GCK(_06648_ ) );
CLKGATE_X1 _14504_ ( .CK(clock ), .E(\u_icache.count_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06649_ ) );
CLKGATE_X1 _14505_ ( .CK(clock ), .E(\u_icache.count_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_06650_ ) );
CLKGATE_X1 _14506_ ( .CK(clock ), .E(\u_icache.count_$_ORNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06651_ ) );
CLKGATE_X1 _14507_ ( .CK(clock ), .E(\u_icache.count_$_OR__B_2_Y_$_ANDNOT__B_Y ), .GCK(_06652_ ) );
CLKGATE_X1 _14508_ ( .CK(clock ), .E(\u_icache.count_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06653_ ) );
CLKGATE_X1 _14509_ ( .CK(clock ), .E(\u_icache.count_$_OR__B_1_Y_$_ANDNOT__B_Y ), .GCK(_06654_ ) );
CLKGATE_X1 _14510_ ( .CK(clock ), .E(icah_ready ), .GCK(_06655_ ) );
CLKGATE_X1 _14511_ ( .CK(clock ), .E(\u_icache.caddr_$_SDFFE_PP0P__Q_E ), .GCK(_06656_ ) );
CLKGATE_X1 _14512_ ( .CK(clock ), .E(\u_exu.exe_start_$_SDFFE_PP0P__Q_E ), .GCK(_06657_ ) );
CLKGATE_X1 _14513_ ( .CK(clock ), .E(\u_exu.exe_end_$_SDFFE_PP0P__Q_E ), .GCK(_06658_ ) );
CLKGATE_X1 _14514_ ( .CK(clock ), .E(\u_exu.alu_p2_$_SDFFE_PP0P__Q_E ), .GCK(_06659_ ) );
CLKGATE_X1 _14515_ ( .CK(clock ), .E(\u_exu.exe_end_$_ANDNOT__B_Y ), .GCK(_06660_ ) );
CLKGATE_X1 _14516_ ( .CK(clock ), .E(flush_$_OR__Y_B ), .GCK(_06661_ ) );
CLKGATE_X1 _14517_ ( .CK(clock ), .E(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_06662_ ) );
CLKGATE_X1 _14518_ ( .CK(clock ), .E(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y ), .GCK(_06663_ ) );
CLKGATE_X1 _14519_ ( .CK(clock ), .E(\u_csr.csr[3]_$_ANDNOT__A_B_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A_$_XOR__A_B_$_OR__A_Y_$_OR__B_1_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_06664_ ) );
CLKGATE_X1 _14520_ ( .CK(clock ), .E(\u_arbiter.wvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06665_ ) );
CLKGATE_X1 _14521_ ( .CK(clock ), .E(\u_arbiter.working_$_SDFFE_PP0P__Q_E ), .GCK(_06666_ ) );
CLKGATE_X1 _14522_ ( .CK(clock ), .E(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_06667_ ) );
CLKGATE_X1 _14523_ ( .CK(clock ), .E(\u_arbiter.rvalid_$_SDFFE_PP0P__Q_E ), .GCK(_06668_ ) );
CLKGATE_X1 _14524_ ( .CK(clock ), .E(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_AND__A_Y ), .GCK(_06669_ ) );
LOGIC1_X1 _14525_ ( .Z(io_master_bready ) );
LOGIC0_X1 _14526_ ( .Z(\io_master_arburst [0] ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q ( .D(_00001_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [31] ), .QN(_07317_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_1 ( .D(_00002_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [30] ), .QN(_07316_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_10 ( .D(_00003_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [21] ), .QN(_07315_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_11 ( .D(_00004_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [20] ), .QN(_07314_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_12 ( .D(_00005_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [19] ), .QN(_07313_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_13 ( .D(_00006_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [18] ), .QN(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_A ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_14 ( .D(_00007_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [17] ), .QN(_07312_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_15 ( .D(_00008_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [16] ), .QN(_07311_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_16 ( .D(_00009_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [15] ), .QN(_07310_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_17 ( .D(_00010_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [14] ), .QN(_07309_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_18 ( .D(_00011_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [13] ), .QN(_07308_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_19 ( .D(_00012_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [12] ), .QN(_07307_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_2 ( .D(_00013_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [29] ), .QN(_07306_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_20 ( .D(_00014_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [11] ), .QN(_07305_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_21 ( .D(_00015_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [10] ), .QN(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_A ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_22 ( .D(_00016_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [9] ), .QN(_07304_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_23 ( .D(_00017_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [8] ), .QN(\u_icache.caddr_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_MUX__B_A ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_24 ( .D(_00018_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [7] ), .QN(_07303_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_25 ( .D(_00019_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [6] ), .QN(\u_icache.caddr_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_MUX__B_A ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_26 ( .D(_00020_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [5] ), .QN(_07302_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_27 ( .D(_00021_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [4] ), .QN(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_A ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_28 ( .D(_00022_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [3] ), .QN(_07301_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_29 ( .D(_00023_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [2] ), .QN(\u_icache.caddr_$_SDFFE_PP0P__Q_29_D_$_MUX__B_A ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_3 ( .D(_00024_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [28] ), .QN(_07300_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_30 ( .D(_00025_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [1] ), .QN(_07299_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_31 ( .D(_00026_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [0] ), .QN(_07298_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_4 ( .D(_00027_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [27] ), .QN(_07297_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_5 ( .D(_00028_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [26] ), .QN(io_master_araddr_$_NOT__Y_5_A_$_MUX__Y_A ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_6 ( .D(_00029_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [25] ), .QN(_07296_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_7 ( .D(_00030_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [24] ), .QN(_07295_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_8 ( .D(_00031_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [23] ), .QN(_07294_ ) );
DFF_X1 \u_arbiter.raddr_$_SDFFE_PP0P__Q_9 ( .D(_00032_ ), .CK(_06669_ ), .Q(\u_arbiter.raddr [22] ), .QN(_07293_ ) );
DFF_X1 \u_arbiter.rmask_$_SDFFE_PP0P__Q ( .D(_00033_ ), .CK(_06669_ ), .Q(\u_arbiter.rmask [1] ), .QN(_07292_ ) );
DFF_X1 \u_arbiter.rmask_$_SDFFE_PP0P__Q_1 ( .D(_00034_ ), .CK(_06669_ ), .Q(\u_arbiter.rmask [0] ), .QN(_07291_ ) );
DFF_X1 \u_arbiter.rsign_$_SDFFE_PP0P__Q ( .D(_00035_ ), .CK(_06669_ ), .Q(\u_arbiter.rsign ), .QN(_07290_ ) );
DFF_X1 \u_arbiter.rvalid_$_SDFFE_PP0P__Q ( .D(_00036_ ), .CK(_06668_ ), .Q(\u_arbiter.rvalid ), .QN(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_A ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q ( .D(_00001_ ), .CK(_06667_ ), .Q(\io_master_awaddr [31] ), .QN(_07289_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_1 ( .D(_00002_ ), .CK(_06667_ ), .Q(\io_master_awaddr [30] ), .QN(_07288_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_10 ( .D(_00003_ ), .CK(_06667_ ), .Q(\io_master_awaddr [21] ), .QN(_07287_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_11 ( .D(_00004_ ), .CK(_06667_ ), .Q(\io_master_awaddr [20] ), .QN(_07286_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_12 ( .D(_00005_ ), .CK(_06667_ ), .Q(\io_master_awaddr [19] ), .QN(_07285_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_13 ( .D(_00006_ ), .CK(_06667_ ), .Q(\io_master_awaddr [18] ), .QN(_07284_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_14 ( .D(_00007_ ), .CK(_06667_ ), .Q(\io_master_awaddr [17] ), .QN(_07283_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_15 ( .D(_00008_ ), .CK(_06667_ ), .Q(\io_master_awaddr [16] ), .QN(_07282_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_16 ( .D(_00009_ ), .CK(_06667_ ), .Q(\io_master_awaddr [15] ), .QN(_07281_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_17 ( .D(_00010_ ), .CK(_06667_ ), .Q(\io_master_awaddr [14] ), .QN(_07280_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_18 ( .D(_00011_ ), .CK(_06667_ ), .Q(\io_master_awaddr [13] ), .QN(_07279_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_19 ( .D(_00012_ ), .CK(_06667_ ), .Q(\io_master_awaddr [12] ), .QN(_07278_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_2 ( .D(_00013_ ), .CK(_06667_ ), .Q(\io_master_awaddr [29] ), .QN(_07277_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_20 ( .D(_00014_ ), .CK(_06667_ ), .Q(\io_master_awaddr [11] ), .QN(_07276_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_21 ( .D(_00015_ ), .CK(_06667_ ), .Q(\io_master_awaddr [10] ), .QN(_07275_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_22 ( .D(_00016_ ), .CK(_06667_ ), .Q(\io_master_awaddr [9] ), .QN(_07274_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_23 ( .D(_00017_ ), .CK(_06667_ ), .Q(\io_master_awaddr [8] ), .QN(_07273_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_24 ( .D(_00018_ ), .CK(_06667_ ), .Q(\io_master_awaddr [7] ), .QN(_07272_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_25 ( .D(_00019_ ), .CK(_06667_ ), .Q(\io_master_awaddr [6] ), .QN(_07271_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_26 ( .D(_00020_ ), .CK(_06667_ ), .Q(\io_master_awaddr [5] ), .QN(_07270_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_27 ( .D(_00021_ ), .CK(_06667_ ), .Q(\io_master_awaddr [4] ), .QN(_07269_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_28 ( .D(_00022_ ), .CK(_06667_ ), .Q(\io_master_awaddr [3] ), .QN(_07268_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_29 ( .D(_00023_ ), .CK(_06667_ ), .Q(\io_master_awaddr [2] ), .QN(_07267_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_3 ( .D(_00024_ ), .CK(_06667_ ), .Q(\io_master_awaddr [28] ), .QN(_07266_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_30 ( .D(_00025_ ), .CK(_06667_ ), .Q(\io_master_awaddr [1] ), .QN(_07265_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_31 ( .D(_00026_ ), .CK(_06667_ ), .Q(\io_master_awaddr [0] ), .QN(_07264_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_4 ( .D(_00027_ ), .CK(_06667_ ), .Q(\io_master_awaddr [27] ), .QN(_07263_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_5 ( .D(_00028_ ), .CK(_06667_ ), .Q(\io_master_awaddr [26] ), .QN(_07262_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_6 ( .D(_00029_ ), .CK(_06667_ ), .Q(\io_master_awaddr [25] ), .QN(_07261_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_7 ( .D(_00030_ ), .CK(_06667_ ), .Q(\io_master_awaddr [24] ), .QN(_07260_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_8 ( .D(_00031_ ), .CK(_06667_ ), .Q(\io_master_awaddr [23] ), .QN(_07259_ ) );
DFF_X1 \u_arbiter.waddr_$_SDFFE_PP0P__Q_9 ( .D(_00032_ ), .CK(_06667_ ), .Q(\io_master_awaddr [22] ), .QN(_07258_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q ( .D(_00037_ ), .CK(_06669_ ), .Q(\u_arbiter.wbaddr [3] ), .QN(_07257_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q_1 ( .D(_00038_ ), .CK(_06669_ ), .Q(\u_arbiter.wbaddr [2] ), .QN(_07256_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q_2 ( .D(_00039_ ), .CK(_06669_ ), .Q(\u_arbiter.wbaddr [1] ), .QN(_07255_ ) );
DFF_X1 \u_arbiter.wbaddr_$_SDFFE_PP0P__Q_3 ( .D(_00040_ ), .CK(_06669_ ), .Q(\u_arbiter.wbaddr [0] ), .QN(_07254_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q ( .D(_00041_ ), .CK(_06667_ ), .Q(\al_wdata [31] ), .QN(_07253_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_1 ( .D(_00042_ ), .CK(_06667_ ), .Q(\al_wdata [30] ), .QN(_07252_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_10 ( .D(_00043_ ), .CK(_06667_ ), .Q(\al_wdata [21] ), .QN(_07251_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_11 ( .D(_00044_ ), .CK(_06667_ ), .Q(\al_wdata [20] ), .QN(_07250_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_12 ( .D(_00045_ ), .CK(_06667_ ), .Q(\al_wdata [19] ), .QN(_07249_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_13 ( .D(_00046_ ), .CK(_06667_ ), .Q(\al_wdata [18] ), .QN(_07248_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_14 ( .D(_00047_ ), .CK(_06667_ ), .Q(\al_wdata [17] ), .QN(_07247_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_15 ( .D(_00048_ ), .CK(_06667_ ), .Q(\al_wdata [16] ), .QN(_07246_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_16 ( .D(_00049_ ), .CK(_06667_ ), .Q(\al_wdata [15] ), .QN(_07245_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_17 ( .D(_00050_ ), .CK(_06667_ ), .Q(\al_wdata [14] ), .QN(_07244_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_18 ( .D(_00051_ ), .CK(_06667_ ), .Q(\al_wdata [13] ), .QN(_07243_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_19 ( .D(_00052_ ), .CK(_06667_ ), .Q(\al_wdata [12] ), .QN(_07242_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_2 ( .D(_00053_ ), .CK(_06667_ ), .Q(\al_wdata [29] ), .QN(_07241_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_20 ( .D(_00054_ ), .CK(_06667_ ), .Q(\al_wdata [11] ), .QN(_07240_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_21 ( .D(_00055_ ), .CK(_06667_ ), .Q(\al_wdata [10] ), .QN(_07239_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_22 ( .D(_00056_ ), .CK(_06667_ ), .Q(\al_wdata [9] ), .QN(_07238_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_23 ( .D(_00057_ ), .CK(_06667_ ), .Q(\al_wdata [8] ), .QN(_07237_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_24 ( .D(_00058_ ), .CK(_06667_ ), .Q(\al_wdata [7] ), .QN(_07236_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_25 ( .D(_00059_ ), .CK(_06667_ ), .Q(\al_wdata [6] ), .QN(_07235_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_26 ( .D(_00060_ ), .CK(_06667_ ), .Q(\al_wdata [5] ), .QN(_07234_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_27 ( .D(_00061_ ), .CK(_06667_ ), .Q(\al_wdata [4] ), .QN(_07233_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_28 ( .D(_00062_ ), .CK(_06667_ ), .Q(\al_wdata [3] ), .QN(_07232_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_29 ( .D(_00063_ ), .CK(_06667_ ), .Q(\al_wdata [2] ), .QN(_07231_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_3 ( .D(_00064_ ), .CK(_06667_ ), .Q(\al_wdata [28] ), .QN(_07230_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_30 ( .D(_00065_ ), .CK(_06667_ ), .Q(\al_wdata [1] ), .QN(_07229_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_31 ( .D(_00066_ ), .CK(_06667_ ), .Q(\al_wdata [0] ), .QN(_07228_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_4 ( .D(_00067_ ), .CK(_06667_ ), .Q(\al_wdata [27] ), .QN(_07227_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_5 ( .D(_00068_ ), .CK(_06667_ ), .Q(\al_wdata [26] ), .QN(_07226_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_6 ( .D(_00069_ ), .CK(_06667_ ), .Q(\al_wdata [25] ), .QN(_07225_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_7 ( .D(_00070_ ), .CK(_06667_ ), .Q(\al_wdata [24] ), .QN(_07224_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_8 ( .D(_00071_ ), .CK(_06667_ ), .Q(\al_wdata [23] ), .QN(_07223_ ) );
DFF_X1 \u_arbiter.wdata_$_SDFFE_PP0P__Q_9 ( .D(_00072_ ), .CK(_06667_ ), .Q(\al_wdata [22] ), .QN(_07222_ ) );
DFF_X1 \u_arbiter.wmask_$_SDFFE_PP0P__Q ( .D(_00033_ ), .CK(_06667_ ), .Q(\al_wmask [1] ), .QN(_07221_ ) );
DFF_X1 \u_arbiter.wmask_$_SDFFE_PP0P__Q_1 ( .D(_00034_ ), .CK(_06667_ ), .Q(\al_wmask [0] ), .QN(_07220_ ) );
DFF_X1 \u_arbiter.working_$_SDFFE_PP0P__Q ( .D(_00073_ ), .CK(_06666_ ), .Q(\u_arbiter.working ), .QN(_07219_ ) );
DFF_X1 \u_arbiter.wvalid_$_SDFFE_PP0P__Q ( .D(_00074_ ), .CK(_06665_ ), .Q(\u_arbiter.wvalid ), .QN(_07218_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q ( .D(_00075_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][31] ), .QN(_07217_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_1 ( .D(_00076_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][30] ), .QN(_07216_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_10 ( .D(_00077_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][21] ), .QN(_07215_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_11 ( .D(_00078_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][20] ), .QN(_07214_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_12 ( .D(_00079_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][19] ), .QN(_07213_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_13 ( .D(_00080_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][18] ), .QN(_07212_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_14 ( .D(_00081_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][17] ), .QN(_07211_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_15 ( .D(_00082_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][16] ), .QN(_07210_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_16 ( .D(_00083_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][15] ), .QN(_07209_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_17 ( .D(_00084_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][14] ), .QN(_07208_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_18 ( .D(_00085_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][13] ), .QN(_07207_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_19 ( .D(_00086_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][10] ), .QN(_07206_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_2 ( .D(_00087_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][29] ), .QN(_07205_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_20 ( .D(_00088_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][9] ), .QN(_07204_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_21 ( .D(_00089_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][8] ), .QN(_07203_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_22 ( .D(_00090_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][7] ), .QN(_07202_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_23 ( .D(_00091_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][6] ), .QN(_07201_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_24 ( .D(_00092_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][5] ), .QN(_07200_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_25 ( .D(_00093_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][4] ), .QN(_07199_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_26 ( .D(_00094_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][3] ), .QN(_07198_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_27 ( .D(_00095_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][2] ), .QN(_07197_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_28 ( .D(_00096_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][1] ), .QN(_07196_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_29 ( .D(_00097_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][0] ), .QN(_07195_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_3 ( .D(_00098_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][28] ), .QN(_07194_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_4 ( .D(_00099_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][27] ), .QN(_07193_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_5 ( .D(_00100_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][26] ), .QN(_07192_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_6 ( .D(_00101_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][25] ), .QN(_07191_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_7 ( .D(_00102_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][24] ), .QN(_07190_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_8 ( .D(_00103_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][23] ), .QN(_07189_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP0P__Q_9 ( .D(_00104_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][22] ), .QN(_07188_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP1P__Q ( .D(_00105_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][12] ), .QN(_07187_ ) );
DFF_X1 \u_csr.csr[0]_$_SDFFE_PP1P__Q_1 ( .D(_00106_ ), .CK(_06664_ ), .Q(\u_csr.csr[0][11] ), .QN(_07186_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q ( .D(_00075_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][31] ), .QN(_07185_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_1 ( .D(_00076_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][30] ), .QN(_07184_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_10 ( .D(_00077_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][21] ), .QN(_07183_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_11 ( .D(_00078_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][20] ), .QN(_07182_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_12 ( .D(_00079_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][19] ), .QN(_07181_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_13 ( .D(_00080_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][18] ), .QN(_07180_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_14 ( .D(_00081_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][17] ), .QN(_07179_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_15 ( .D(_00082_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][16] ), .QN(_07178_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_16 ( .D(_00083_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][15] ), .QN(_07177_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_17 ( .D(_00084_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][14] ), .QN(_07176_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_18 ( .D(_00085_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][13] ), .QN(_07175_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_19 ( .D(_00107_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][12] ), .QN(_07174_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_2 ( .D(_00087_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][29] ), .QN(_07173_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_20 ( .D(_00108_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][11] ), .QN(_07172_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_21 ( .D(_00086_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][10] ), .QN(_07171_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_22 ( .D(_00088_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][9] ), .QN(_07170_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_23 ( .D(_00089_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][8] ), .QN(_07169_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_24 ( .D(_00090_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][7] ), .QN(_07168_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_25 ( .D(_00091_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][6] ), .QN(_07167_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_26 ( .D(_00092_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][5] ), .QN(_07166_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_27 ( .D(_00093_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][4] ), .QN(_07165_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_28 ( .D(_00094_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][3] ), .QN(_07164_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_29 ( .D(_00095_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][2] ), .QN(_07163_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_3 ( .D(_00098_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][28] ), .QN(_07162_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_30 ( .D(_00096_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][1] ), .QN(_07161_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_31 ( .D(_00097_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][0] ), .QN(_07160_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_4 ( .D(_00099_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][27] ), .QN(_07159_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_5 ( .D(_00100_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][26] ), .QN(_07158_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_6 ( .D(_00101_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][25] ), .QN(_07157_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_7 ( .D(_00102_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][24] ), .QN(_07156_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_8 ( .D(_00103_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][23] ), .QN(_07155_ ) );
DFF_X1 \u_csr.csr[1]_$_SDFFE_PP0P__Q_9 ( .D(_00104_ ), .CK(_06663_ ), .Q(\u_csr.csr[1][22] ), .QN(_07154_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q ( .D(_00075_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][31] ), .QN(_07153_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_1 ( .D(_00076_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][30] ), .QN(_07152_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_10 ( .D(_00077_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][21] ), .QN(_07151_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_11 ( .D(_00078_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][20] ), .QN(_07150_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_12 ( .D(_00079_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][19] ), .QN(_07149_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_13 ( .D(_00080_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][18] ), .QN(_07148_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_14 ( .D(_00081_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][17] ), .QN(_07147_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_15 ( .D(_00082_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][16] ), .QN(_07146_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_16 ( .D(_00083_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][15] ), .QN(_07145_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_17 ( .D(_00084_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][14] ), .QN(_07144_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_18 ( .D(_00085_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][13] ), .QN(_07143_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_19 ( .D(_00107_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][12] ), .QN(_07142_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_2 ( .D(_00087_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][29] ), .QN(_07141_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_20 ( .D(_00108_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][11] ), .QN(_07140_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_21 ( .D(_00086_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][10] ), .QN(_07139_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_22 ( .D(_00088_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][9] ), .QN(_07138_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_23 ( .D(_00089_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][8] ), .QN(_07137_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_24 ( .D(_00090_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][7] ), .QN(_07136_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_25 ( .D(_00091_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][6] ), .QN(_07135_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_26 ( .D(_00092_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][5] ), .QN(_07134_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_27 ( .D(_00093_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][4] ), .QN(_07133_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_28 ( .D(_00094_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][3] ), .QN(_07132_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_29 ( .D(_00095_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][2] ), .QN(_07131_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_3 ( .D(_00098_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][28] ), .QN(_07130_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_30 ( .D(_00096_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][1] ), .QN(_07129_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_31 ( .D(_00097_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][0] ), .QN(_07128_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_4 ( .D(_00099_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][27] ), .QN(_07127_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_5 ( .D(_00100_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][26] ), .QN(_07126_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_6 ( .D(_00101_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][25] ), .QN(_07125_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_7 ( .D(_00102_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][24] ), .QN(_07124_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_8 ( .D(_00103_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][23] ), .QN(_07123_ ) );
DFF_X1 \u_csr.csr[2]_$_SDFFE_PP0P__Q_9 ( .D(_00104_ ), .CK(_06662_ ), .Q(\u_csr.csr[2][22] ), .QN(_07122_ ) );
DFF_X1 \u_csr.csr[3]_$_SDFFCE_PN0P__Q ( .D(_00109_ ), .CK(_06661_ ), .Q(\u_csr.csr[3][0] ), .QN(_07121_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q ( .D(_00110_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [11] ), .QN(_07120_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_1 ( .D(_00111_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [10] ), .QN(_07119_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_10 ( .D(_00112_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [1] ), .QN(_07118_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_11 ( .D(_00113_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [0] ), .QN(_07117_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_2 ( .D(_00114_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [9] ), .QN(_07116_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_3 ( .D(_00115_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [8] ), .QN(_07115_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_4 ( .D(_00116_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [7] ), .QN(_07114_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_5 ( .D(_00117_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [6] ), .QN(_07113_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_6 ( .D(_00118_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [5] ), .QN(_07112_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_7 ( .D(_00119_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [4] ), .QN(_07111_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_8 ( .D(_00120_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [3] ), .QN(_07110_ ) );
DFF_X1 \u_exu.acsrd_$_SDFFE_PP0P__Q_9 ( .D(_00121_ ), .CK(_06660_ ), .Q(\u_exu.acsrd [2] ), .QN(_07109_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q ( .D(_00122_ ), .CK(_06659_ ), .Q(\u_exu.alu_ctrl [6] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_1 ( .D(_00123_ ), .CK(_06659_ ), .Q(\u_exu.alu_ctrl [5] ), .QN(_07108_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_2 ( .D(_00124_ ), .CK(_06659_ ), .Q(\u_exu.alu_ctrl [4] ), .QN(_07107_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_3 ( .D(_00125_ ), .CK(_06659_ ), .Q(\u_exu.alu_ctrl [3] ), .QN(_07106_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_4 ( .D(_00126_ ), .CK(_06659_ ), .Q(\u_exu.alu_ctrl [2] ), .QN(_07105_ ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_5 ( .D(_00127_ ), .CK(_06659_ ), .Q(\u_exu.alu_ctrl [1] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_Y_$_MUX__B_A_$_NOR__Y_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_exu.alu_ctrl_$_SDFFE_PP0P__Q_6 ( .D(_00128_ ), .CK(_06659_ ), .Q(\u_exu.alu_ctrl [0] ), .QN(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q ( .D(_00129_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [31] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_1 ( .D(_00130_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [30] ), .QN(_07104_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_10 ( .D(_00131_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [21] ), .QN(\u_exu.rd_$_MUX__Y_9_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_11 ( .D(_00132_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [20] ), .QN(_07103_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_12 ( .D(_00133_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [19] ), .QN(\u_exu.rd_$_MUX__Y_12_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_13 ( .D(_00134_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [18] ), .QN(_07102_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_14 ( .D(_00135_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [17] ), .QN(\u_exu.rd_$_MUX__Y_13_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_15 ( .D(_00136_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [16] ), .QN(_07101_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_16 ( .D(_00137_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [15] ), .QN(\u_exu.rd_$_MUX__Y_16_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_17 ( .D(_00138_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [14] ), .QN(_07100_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_18 ( .D(_00139_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [13] ), .QN(_07099_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_19 ( .D(_00140_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [12] ), .QN(_07098_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_2 ( .D(_00141_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [29] ), .QN(_07097_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_20 ( .D(_00142_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [11] ), .QN(\u_exu.rd_$_MUX__Y_20_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_21 ( .D(_00143_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [10] ), .QN(_07096_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_22 ( .D(_00144_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [9] ), .QN(\u_exu.rd_$_MUX__Y_21_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_23 ( .D(_00145_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [8] ), .QN(_07095_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_24 ( .D(_00146_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [7] ), .QN(\u_exu.rd_$_MUX__Y_24_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_25 ( .D(_00147_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [6] ), .QN(_07094_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_26 ( .D(_00148_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [5] ), .QN(\u_exu.rd_$_MUX__Y_25_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_27 ( .D(_00149_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [4] ), .QN(_07093_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_28 ( .D(_00150_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [3] ), .QN(\u_exu.rd_$_MUX__Y_28_A_$_MUX__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_29 ( .D(_00151_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [2] ), .QN(_07092_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_3 ( .D(_00152_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [28] ), .QN(_07091_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_30 ( .D(_00153_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [1] ), .QN(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_31 ( .D(_00154_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [0] ), .QN(\u_exu.rd_$_MUX__Y_30_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_4 ( .D(_00155_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [27] ), .QN(_07090_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_5 ( .D(_00156_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [26] ), .QN(_07089_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_6 ( .D(_00157_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [25] ), .QN(_07088_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_7 ( .D(_00158_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [24] ), .QN(_07087_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_8 ( .D(_00159_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [23] ), .QN(_07086_ ) );
DFF_X1 \u_exu.alu_p1_$_SDFFE_PP0P__Q_9 ( .D(_00160_ ), .CK(_06659_ ), .Q(\u_exu.alu_p1 [22] ), .QN(_07085_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q ( .D(_00161_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [31] ), .QN(_07084_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_1 ( .D(_00162_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [30] ), .QN(_07083_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_10 ( .D(_00163_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [21] ), .QN(_07082_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_11 ( .D(_00164_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [20] ), .QN(_07081_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_12 ( .D(_00165_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [19] ), .QN(_07080_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_13 ( .D(_00166_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [18] ), .QN(_07079_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_14 ( .D(_00167_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [17] ), .QN(_07078_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_15 ( .D(_00168_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [16] ), .QN(_07077_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_16 ( .D(_00169_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [15] ), .QN(_07076_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_17 ( .D(_00170_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [14] ), .QN(_07075_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_18 ( .D(_00171_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [13] ), .QN(_07074_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_19 ( .D(_00172_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [12] ), .QN(_07073_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_2 ( .D(_00173_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [29] ), .QN(_07072_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_20 ( .D(_00174_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [11] ), .QN(_07071_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_21 ( .D(_00175_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [10] ), .QN(_07070_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_22 ( .D(_00176_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [9] ), .QN(_07069_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_23 ( .D(_00177_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [8] ), .QN(_07068_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_24 ( .D(_00178_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [7] ), .QN(_07067_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_25 ( .D(_00179_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [6] ), .QN(_07066_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_26 ( .D(_00180_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [5] ), .QN(_07065_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_27 ( .D(_00181_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [4] ), .QN(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_B_$_MUX__B_A_$_NAND__Y_B ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_28 ( .D(_00182_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [3] ), .QN(_07064_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_29 ( .D(_00183_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [2] ), .QN(_07063_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_3 ( .D(_00184_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [28] ), .QN(_07062_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_30 ( .D(_00185_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [1] ), .QN(_07061_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_31 ( .D(_00186_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [0] ), .QN(_07060_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_4 ( .D(_00187_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [27] ), .QN(_07059_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_5 ( .D(_00188_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [26] ), .QN(_07058_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_6 ( .D(_00189_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [25] ), .QN(_07057_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_7 ( .D(_00190_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [24] ), .QN(_07056_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_8 ( .D(_00191_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [23] ), .QN(_07055_ ) );
DFF_X1 \u_exu.alu_p2_$_SDFFE_PP0P__Q_9 ( .D(_00192_ ), .CK(_06659_ ), .Q(\u_exu.alu_p2 [22] ), .QN(_07054_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q ( .D(_00193_ ), .CK(_06660_ ), .Q(\ea_ard [3] ), .QN(_07053_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q_1 ( .D(_00194_ ), .CK(_06660_ ), .Q(\ea_ard [2] ), .QN(_07052_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q_2 ( .D(_00195_ ), .CK(_06660_ ), .Q(\ea_ard [1] ), .QN(_07051_ ) );
DFF_X1 \u_exu.ard_$_SDFFE_PP0P__Q_3 ( .D(_00196_ ), .CK(_06660_ ), .Q(\ea_ard [0] ), .QN(_07050_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q ( .D(_00197_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [31] ), .QN(_07049_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_1 ( .D(_00198_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [30] ), .QN(_07048_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_10 ( .D(_00199_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [21] ), .QN(_07047_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_11 ( .D(_00200_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [20] ), .QN(_07046_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_12 ( .D(_00201_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [19] ), .QN(_07045_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_13 ( .D(_00202_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [18] ), .QN(_07044_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_14 ( .D(_00203_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [17] ), .QN(_07043_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_15 ( .D(_00204_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [16] ), .QN(_07042_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_16 ( .D(_00205_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [15] ), .QN(_07041_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_17 ( .D(_00206_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [14] ), .QN(_07040_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_18 ( .D(_00207_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [13] ), .QN(_07039_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_19 ( .D(_00208_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [12] ), .QN(_07038_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_2 ( .D(_00209_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [29] ), .QN(_07037_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_20 ( .D(_00210_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [11] ), .QN(_07036_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_21 ( .D(_00211_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [10] ), .QN(_07035_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_22 ( .D(_00212_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [9] ), .QN(_07034_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_23 ( .D(_00213_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [8] ), .QN(_07033_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_24 ( .D(_00214_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [7] ), .QN(_07032_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_25 ( .D(_00215_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [6] ), .QN(_07031_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_26 ( .D(_00216_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [5] ), .QN(_07030_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_27 ( .D(_00217_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [4] ), .QN(_07029_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_28 ( .D(_00218_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [3] ), .QN(_07028_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_29 ( .D(_00219_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [2] ), .QN(_07027_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_3 ( .D(_00220_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [28] ), .QN(_07026_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_30 ( .D(_00221_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [1] ), .QN(_07025_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_31 ( .D(_00222_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [0] ), .QN(_07024_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_4 ( .D(_00223_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [27] ), .QN(_07023_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_5 ( .D(_00224_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [26] ), .QN(_07022_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_6 ( .D(_00225_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [25] ), .QN(_07021_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_7 ( .D(_00226_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [24] ), .QN(_07020_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_8 ( .D(_00227_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [23] ), .QN(_07019_ ) );
DFF_X1 \u_exu.ecsr_$_SDFFE_PP0P__Q_9 ( .D(_00228_ ), .CK(_06660_ ), .Q(\u_exu.ecsr [22] ), .QN(_07018_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q ( .D(_00229_ ), .CK(_06660_ ), .Q(\u_exu.eopt [15] ), .QN(_07017_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_1 ( .D(_00230_ ), .CK(_06660_ ), .Q(ea_rsign ), .QN(_07016_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_2 ( .D(_00231_ ), .CK(_06660_ ), .Q(\u_exu.eopt [12] ), .QN(_07015_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_3 ( .D(_00232_ ), .CK(_06660_ ), .Q(\ea_mask [1] ), .QN(_07014_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_4 ( .D(_00233_ ), .CK(_06660_ ), .Q(\ea_mask [0] ), .QN(_07013_ ) );
DFF_X1 \u_exu.eopt_$_SDFFE_PP0P__Q_5 ( .D(_00234_ ), .CK(_06660_ ), .Q(\u_exu.eopt [0] ), .QN(_07012_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q ( .D(_00235_ ), .CK(_06660_ ), .Q(\ea_pc [31] ), .QN(_07011_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_1 ( .D(_00236_ ), .CK(_06660_ ), .Q(\ea_pc [30] ), .QN(_07010_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_10 ( .D(_00237_ ), .CK(_06660_ ), .Q(\ea_pc [21] ), .QN(_07009_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_11 ( .D(_00238_ ), .CK(_06660_ ), .Q(\ea_pc [20] ), .QN(_07008_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_12 ( .D(_00239_ ), .CK(_06660_ ), .Q(\ea_pc [19] ), .QN(_07007_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_13 ( .D(_00240_ ), .CK(_06660_ ), .Q(\ea_pc [18] ), .QN(_07006_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_14 ( .D(_00241_ ), .CK(_06660_ ), .Q(\ea_pc [17] ), .QN(_07005_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_15 ( .D(_00242_ ), .CK(_06660_ ), .Q(\ea_pc [16] ), .QN(_07004_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_16 ( .D(_00243_ ), .CK(_06660_ ), .Q(\ea_pc [15] ), .QN(_07003_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_17 ( .D(_00244_ ), .CK(_06660_ ), .Q(\ea_pc [14] ), .QN(_07002_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_18 ( .D(_00245_ ), .CK(_06660_ ), .Q(\ea_pc [13] ), .QN(_07001_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_19 ( .D(_00246_ ), .CK(_06660_ ), .Q(\ea_pc [12] ), .QN(_07000_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_2 ( .D(_00247_ ), .CK(_06660_ ), .Q(\ea_pc [29] ), .QN(_06999_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_20 ( .D(_00248_ ), .CK(_06660_ ), .Q(\ea_pc [11] ), .QN(_06998_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_21 ( .D(_00249_ ), .CK(_06660_ ), .Q(\ea_pc [10] ), .QN(_06997_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_22 ( .D(_00250_ ), .CK(_06660_ ), .Q(\ea_pc [9] ), .QN(_06996_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_23 ( .D(_00251_ ), .CK(_06660_ ), .Q(\ea_pc [8] ), .QN(_06995_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_24 ( .D(_00252_ ), .CK(_06660_ ), .Q(\ea_pc [7] ), .QN(_06994_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_25 ( .D(_00253_ ), .CK(_06660_ ), .Q(\ea_pc [6] ), .QN(_06993_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_26 ( .D(_00254_ ), .CK(_06660_ ), .Q(\ea_pc [5] ), .QN(_06992_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_27 ( .D(_00255_ ), .CK(_06660_ ), .Q(\ea_pc [4] ), .QN(_06991_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_28 ( .D(_00256_ ), .CK(_06660_ ), .Q(\ea_pc [3] ), .QN(_06990_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_29 ( .D(_00257_ ), .CK(_06660_ ), .Q(\ea_pc [2] ), .QN(_06989_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_3 ( .D(_00258_ ), .CK(_06660_ ), .Q(\ea_pc [28] ), .QN(_06988_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_30 ( .D(_00259_ ), .CK(_06660_ ), .Q(\ea_pc [1] ), .QN(_06987_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_31 ( .D(_00260_ ), .CK(_06660_ ), .Q(\ea_pc [0] ), .QN(_06986_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_4 ( .D(_00261_ ), .CK(_06660_ ), .Q(\ea_pc [27] ), .QN(_06985_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_5 ( .D(_00262_ ), .CK(_06660_ ), .Q(\ea_pc [26] ), .QN(_06984_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_6 ( .D(_00263_ ), .CK(_06660_ ), .Q(\ea_pc [25] ), .QN(_06983_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_7 ( .D(_00264_ ), .CK(_06660_ ), .Q(\ea_pc [24] ), .QN(_06982_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_8 ( .D(_00265_ ), .CK(_06660_ ), .Q(\ea_pc [23] ), .QN(_06981_ ) );
DFF_X1 \u_exu.epc_$_SDFFE_PP0P__Q_9 ( .D(_00266_ ), .CK(_06660_ ), .Q(\ea_pc [22] ), .QN(_06980_ ) );
DFF_X1 \u_exu.error_$_SDFFE_PP0P__Q ( .D(_00267_ ), .CK(_06660_ ), .Q(ea_err ), .QN(\u_arbiter.working_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__B_A ) );
DFF_X1 \u_exu.errtp_$_SDFFE_PP0P__Q ( .D(_00268_ ), .CK(_06660_ ), .Q(\ea_errtp [0] ), .QN(_06979_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q ( .D(_00269_ ), .CK(_06660_ ), .Q(\ea_wdata [31] ), .QN(_06978_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_1 ( .D(_00270_ ), .CK(_06660_ ), .Q(\ea_wdata [30] ), .QN(_06977_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_10 ( .D(_00271_ ), .CK(_06660_ ), .Q(\ea_wdata [21] ), .QN(_06976_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_11 ( .D(_00272_ ), .CK(_06660_ ), .Q(\ea_wdata [20] ), .QN(_06975_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_12 ( .D(_00273_ ), .CK(_06660_ ), .Q(\ea_wdata [19] ), .QN(_06974_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_13 ( .D(_00274_ ), .CK(_06660_ ), .Q(\ea_wdata [18] ), .QN(_06973_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_14 ( .D(_00275_ ), .CK(_06660_ ), .Q(\ea_wdata [17] ), .QN(_06972_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_15 ( .D(_00276_ ), .CK(_06660_ ), .Q(\ea_wdata [16] ), .QN(_06971_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_16 ( .D(_00277_ ), .CK(_06660_ ), .Q(\ea_wdata [15] ), .QN(_06970_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_17 ( .D(_00278_ ), .CK(_06660_ ), .Q(\ea_wdata [14] ), .QN(_06969_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_18 ( .D(_00279_ ), .CK(_06660_ ), .Q(\ea_wdata [13] ), .QN(_06968_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_19 ( .D(_00280_ ), .CK(_06660_ ), .Q(\ea_wdata [12] ), .QN(_06967_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_2 ( .D(_00281_ ), .CK(_06660_ ), .Q(\ea_wdata [29] ), .QN(_06966_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_20 ( .D(_00282_ ), .CK(_06660_ ), .Q(\ea_wdata [11] ), .QN(_06965_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_21 ( .D(_00283_ ), .CK(_06660_ ), .Q(\ea_wdata [10] ), .QN(_06964_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_22 ( .D(_00284_ ), .CK(_06660_ ), .Q(\ea_wdata [9] ), .QN(_06963_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_23 ( .D(_00285_ ), .CK(_06660_ ), .Q(\ea_wdata [8] ), .QN(_06962_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_24 ( .D(_00286_ ), .CK(_06660_ ), .Q(\ea_wdata [7] ), .QN(_06961_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_25 ( .D(_00287_ ), .CK(_06660_ ), .Q(\ea_wdata [6] ), .QN(_06960_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_26 ( .D(_00288_ ), .CK(_06660_ ), .Q(\ea_wdata [5] ), .QN(_06959_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_27 ( .D(_00289_ ), .CK(_06660_ ), .Q(\ea_wdata [4] ), .QN(_06958_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_28 ( .D(_00290_ ), .CK(_06660_ ), .Q(\ea_wdata [3] ), .QN(_06957_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_29 ( .D(_00291_ ), .CK(_06660_ ), .Q(\ea_wdata [2] ), .QN(_06956_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_3 ( .D(_00292_ ), .CK(_06660_ ), .Q(\ea_wdata [28] ), .QN(_06955_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_30 ( .D(_00293_ ), .CK(_06660_ ), .Q(\ea_wdata [1] ), .QN(_06954_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_31 ( .D(_00294_ ), .CK(_06660_ ), .Q(\ea_wdata [0] ), .QN(_06953_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_4 ( .D(_00295_ ), .CK(_06660_ ), .Q(\ea_wdata [27] ), .QN(_06952_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_5 ( .D(_00296_ ), .CK(_06660_ ), .Q(\ea_wdata [26] ), .QN(_06951_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_6 ( .D(_00297_ ), .CK(_06660_ ), .Q(\ea_wdata [25] ), .QN(_06950_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_7 ( .D(_00298_ ), .CK(_06660_ ), .Q(\ea_wdata [24] ), .QN(_06949_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_8 ( .D(_00299_ ), .CK(_06660_ ), .Q(\ea_wdata [23] ), .QN(_06948_ ) );
DFF_X1 \u_exu.ers2_$_SDFFE_PP0P__Q_9 ( .D(_00300_ ), .CK(_06660_ ), .Q(\ea_wdata [22] ), .QN(_06947_ ) );
DFF_X1 \u_exu.exe_end_$_SDFFE_PP0P__Q ( .D(_00301_ ), .CK(_06658_ ), .Q(exu_valid ), .QN(_06946_ ) );
DFF_X1 \u_exu.exe_start_$_SDFFE_PP0P__Q ( .D(_00302_ ), .CK(_06657_ ), .Q(\u_exu.exe_start ), .QN(_06945_ ) );
DFF_X1 \u_exu.jmpc_ok_$_SDFF_PP0__Q ( .D(_00304_ ), .CK(clock ), .Q(\u_exu.jmpc_ok ), .QN(_06943_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q ( .D(_00303_ ), .CK(_06660_ ), .Q(\ea_addr [31] ), .QN(_06944_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_1 ( .D(_00305_ ), .CK(_06660_ ), .Q(\ea_addr [30] ), .QN(_06942_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_10 ( .D(_00306_ ), .CK(_06660_ ), .Q(\ea_addr [21] ), .QN(_06941_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_11 ( .D(_00307_ ), .CK(_06660_ ), .Q(\ea_addr [20] ), .QN(_06940_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_12 ( .D(_00308_ ), .CK(_06660_ ), .Q(\ea_addr [19] ), .QN(_06939_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_13 ( .D(_00309_ ), .CK(_06660_ ), .Q(\ea_addr [18] ), .QN(_06938_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_14 ( .D(_00310_ ), .CK(_06660_ ), .Q(\ea_addr [17] ), .QN(_06937_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_15 ( .D(_00311_ ), .CK(_06660_ ), .Q(\ea_addr [16] ), .QN(_06936_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_16 ( .D(_00312_ ), .CK(_06660_ ), .Q(\ea_addr [15] ), .QN(_06935_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_17 ( .D(_00313_ ), .CK(_06660_ ), .Q(\ea_addr [14] ), .QN(_06934_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_18 ( .D(_00314_ ), .CK(_06660_ ), .Q(\ea_addr [13] ), .QN(_06933_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_19 ( .D(_00315_ ), .CK(_06660_ ), .Q(\ea_addr [12] ), .QN(_06932_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_2 ( .D(_00316_ ), .CK(_06660_ ), .Q(\ea_addr [29] ), .QN(_06931_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_20 ( .D(_00317_ ), .CK(_06660_ ), .Q(\ea_addr [11] ), .QN(_06930_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_21 ( .D(_00318_ ), .CK(_06660_ ), .Q(\ea_addr [10] ), .QN(_06929_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_22 ( .D(_00319_ ), .CK(_06660_ ), .Q(\ea_addr [9] ), .QN(_06928_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_23 ( .D(_00320_ ), .CK(_06660_ ), .Q(\ea_addr [8] ), .QN(_06927_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_24 ( .D(_00321_ ), .CK(_06660_ ), .Q(\ea_addr [7] ), .QN(_06926_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_25 ( .D(_00322_ ), .CK(_06660_ ), .Q(\ea_addr [6] ), .QN(_06925_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_26 ( .D(_00323_ ), .CK(_06660_ ), .Q(\ea_addr [5] ), .QN(_06924_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_27 ( .D(_00324_ ), .CK(_06660_ ), .Q(\ea_addr [4] ), .QN(_06923_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_28 ( .D(_00325_ ), .CK(_06660_ ), .Q(\ea_addr [3] ), .QN(_06922_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_29 ( .D(_00326_ ), .CK(_06660_ ), .Q(\ea_addr [2] ), .QN(_06921_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_3 ( .D(_00327_ ), .CK(_06660_ ), .Q(\ea_addr [28] ), .QN(_06920_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_30 ( .D(_00328_ ), .CK(_06660_ ), .Q(\ea_addr [1] ), .QN(_06919_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_31 ( .D(_00329_ ), .CK(_06660_ ), .Q(\ea_addr [0] ), .QN(_06918_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_4 ( .D(_00330_ ), .CK(_06660_ ), .Q(\ea_addr [27] ), .QN(_06917_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_5 ( .D(_00331_ ), .CK(_06660_ ), .Q(\ea_addr [26] ), .QN(_06916_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_6 ( .D(_00332_ ), .CK(_06660_ ), .Q(\ea_addr [25] ), .QN(_06915_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_7 ( .D(_00333_ ), .CK(_06660_ ), .Q(\ea_addr [24] ), .QN(_06914_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_8 ( .D(_00334_ ), .CK(_06660_ ), .Q(\ea_addr [23] ), .QN(_06913_ ) );
DFF_X1 \u_exu.rdo_$_SDFFE_PP0P__Q_9 ( .D(_00335_ ), .CK(_06660_ ), .Q(\ea_addr [22] ), .QN(_06912_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q ( .D(_00337_ ), .CK(clock ), .Q(\u_exu.rlock [15] ), .QN(_06910_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_1 ( .D(_00338_ ), .CK(clock ), .Q(\u_exu.rlock [14] ), .QN(_06909_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_10 ( .D(_00339_ ), .CK(clock ), .Q(\u_exu.rlock [5] ), .QN(_06908_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_11 ( .D(_00340_ ), .CK(clock ), .Q(\u_exu.rlock [4] ), .QN(_06907_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_12 ( .D(_00341_ ), .CK(clock ), .Q(\u_exu.rlock [3] ), .QN(_06906_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_13 ( .D(_00342_ ), .CK(clock ), .Q(\u_exu.rlock [2] ), .QN(_06905_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_14 ( .D(_00343_ ), .CK(clock ), .Q(\u_exu.rlock [1] ), .QN(_06904_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_15 ( .D(_00344_ ), .CK(clock ), .Q(\u_exu.rlock [0] ), .QN(_06903_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_2 ( .D(_00345_ ), .CK(clock ), .Q(\u_exu.rlock [13] ), .QN(_06902_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_3 ( .D(_00346_ ), .CK(clock ), .Q(\u_exu.rlock [12] ), .QN(_06901_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_4 ( .D(_00347_ ), .CK(clock ), .Q(\u_exu.rlock [11] ), .QN(_06900_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_5 ( .D(_00348_ ), .CK(clock ), .Q(\u_exu.rlock [10] ), .QN(_06899_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_6 ( .D(_00349_ ), .CK(clock ), .Q(\u_exu.rlock [9] ), .QN(_06898_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_7 ( .D(_00350_ ), .CK(clock ), .Q(\u_exu.rlock [8] ), .QN(_06897_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_8 ( .D(_00351_ ), .CK(clock ), .Q(\u_exu.rlock [7] ), .QN(_06896_ ) );
DFF_X1 \u_exu.rlock_$_SDFF_PP0__Q_9 ( .D(_00352_ ), .CK(clock ), .Q(\u_exu.rlock [6] ), .QN(_06895_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q ( .D(_00336_ ), .CK(_06656_ ), .Q(\ca_addr [31] ), .QN(_06911_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_1 ( .D(_00353_ ), .CK(_06656_ ), .Q(\ca_addr [30] ), .QN(_06894_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_10 ( .D(_00354_ ), .CK(_06656_ ), .Q(\ca_addr [21] ), .QN(_06893_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_11 ( .D(_00355_ ), .CK(_06656_ ), .Q(\ca_addr [20] ), .QN(_06892_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_12 ( .D(_00356_ ), .CK(_06656_ ), .Q(\ca_addr [19] ), .QN(_06891_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_13 ( .D(_00357_ ), .CK(_06656_ ), .Q(\ca_addr [18] ), .QN(io_master_araddr_$_NOT__Y_4_A_$_MUX__Y_B ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_14 ( .D(_00358_ ), .CK(_06656_ ), .Q(\ca_addr [17] ), .QN(_06890_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_15 ( .D(_00359_ ), .CK(_06656_ ), .Q(\ca_addr [16] ), .QN(_06889_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_16 ( .D(_00360_ ), .CK(_06656_ ), .Q(\ca_addr [15] ), .QN(_06888_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_17 ( .D(_00361_ ), .CK(_06656_ ), .Q(\ca_addr [14] ), .QN(_06887_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_18 ( .D(_00362_ ), .CK(_06656_ ), .Q(\ca_addr [13] ), .QN(_06886_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_19 ( .D(_00363_ ), .CK(_06656_ ), .Q(\ca_addr [12] ), .QN(_06885_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_2 ( .D(_00364_ ), .CK(_06656_ ), .Q(\ca_addr [29] ), .QN(_06884_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_20 ( .D(_00365_ ), .CK(_06656_ ), .Q(\ca_addr [11] ), .QN(_06883_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_21 ( .D(_00366_ ), .CK(_06656_ ), .Q(\ca_addr [10] ), .QN(io_master_araddr_$_NOT__Y_3_A_$_MUX__Y_B ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_22 ( .D(_00367_ ), .CK(_06656_ ), .Q(\ca_addr [9] ), .QN(_06882_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_23 ( .D(_00368_ ), .CK(_06656_ ), .Q(\ca_addr [8] ), .QN(\u_icache.caddr_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_24 ( .D(_00369_ ), .CK(_06656_ ), .Q(\ca_addr [7] ), .QN(_06881_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_25 ( .D(_00370_ ), .CK(_06656_ ), .Q(\ca_addr [6] ), .QN(\u_icache.caddr_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_26 ( .D(_00371_ ), .CK(_06656_ ), .Q(\ca_addr [5] ), .QN(_06880_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_27 ( .D(_00372_ ), .CK(_06656_ ), .Q(\ca_addr [4] ), .QN(io_master_araddr_$_NOT__Y_2_A_$_MUX__Y_B ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_28 ( .D(_00373_ ), .CK(_06655_ ), .Q(\ca_addr [3] ), .QN(_06879_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_29 ( .D(_00374_ ), .CK(_06655_ ), .Q(\ca_addr [2] ), .QN(\u_icache.caddr_$_SDFFE_PP0P__Q_28_D [0] ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_3 ( .D(_00375_ ), .CK(_06656_ ), .Q(\ca_addr [28] ), .QN(_06878_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_4 ( .D(_00376_ ), .CK(_06656_ ), .Q(\ca_addr [27] ), .QN(_06877_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_5 ( .D(_00377_ ), .CK(_06656_ ), .Q(\ca_addr [26] ), .QN(io_master_araddr_$_NOT__Y_5_A_$_MUX__Y_B ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_6 ( .D(_00378_ ), .CK(_06656_ ), .Q(\ca_addr [25] ), .QN(_06876_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_7 ( .D(_00379_ ), .CK(_06656_ ), .Q(\ca_addr [24] ), .QN(_06875_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_8 ( .D(_00380_ ), .CK(_06656_ ), .Q(\ca_addr [23] ), .QN(_06874_ ) );
DFF_X1 \u_icache.caddr_$_SDFFE_PP0P__Q_9 ( .D(_00381_ ), .CK(_06656_ ), .Q(\ca_addr [22] ), .QN(_07318_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][31] ), .QN(_07319_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][30] ), .QN(_07320_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][21] ), .QN(_07321_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][20] ), .QN(_07322_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][19] ), .QN(_07323_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][18] ), .QN(_07324_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][17] ), .QN(_07325_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][16] ), .QN(_07326_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][15] ), .QN(_07327_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][14] ), .QN(_07328_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][13] ), .QN(_07329_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][12] ), .QN(_07330_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][29] ), .QN(_07331_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][11] ), .QN(_07332_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][10] ), .QN(_07333_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][9] ), .QN(_07334_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][8] ), .QN(_07335_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][7] ), .QN(_07336_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][6] ), .QN(_07337_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][5] ), .QN(_07338_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][4] ), .QN(_07339_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][3] ), .QN(_07340_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][2] ), .QN(_07341_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][28] ), .QN(_07342_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][1] ), .QN(_07343_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][0] ), .QN(_07344_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][27] ), .QN(_07345_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][26] ), .QN(_07346_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][25] ), .QN(_07347_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][24] ), .QN(_07348_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][23] ), .QN(_07349_ ) );
DFF_X1 \u_icache.cblocks[0]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06654_ ), .Q(\u_icache.cblocks[0][22] ), .QN(_07350_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][31] ), .QN(_07351_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][30] ), .QN(_07352_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][21] ), .QN(_07353_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][20] ), .QN(_07354_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][19] ), .QN(_07355_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][18] ), .QN(_07356_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][17] ), .QN(_07357_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][16] ), .QN(_07358_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][15] ), .QN(_07359_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][14] ), .QN(_07360_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][13] ), .QN(_07361_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][12] ), .QN(_07362_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][29] ), .QN(_07363_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][11] ), .QN(_07364_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][10] ), .QN(_07365_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][9] ), .QN(_07366_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][8] ), .QN(_07367_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][7] ), .QN(_07368_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][6] ), .QN(_07369_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][5] ), .QN(_07370_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][4] ), .QN(_07371_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][3] ), .QN(_07372_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][2] ), .QN(_07373_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][28] ), .QN(_07374_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][1] ), .QN(_07375_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][0] ), .QN(_07376_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][27] ), .QN(_07377_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][26] ), .QN(_07378_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][25] ), .QN(_07379_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][24] ), .QN(_07380_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][23] ), .QN(_07381_ ) );
DFF_X1 \u_icache.cblocks[1]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06653_ ), .Q(\u_icache.cblocks[1][22] ), .QN(_07382_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][31] ), .QN(_07383_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][30] ), .QN(_07384_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][21] ), .QN(_07385_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][20] ), .QN(_07386_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][19] ), .QN(_07387_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][18] ), .QN(_07388_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][17] ), .QN(_07389_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][16] ), .QN(_07390_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][15] ), .QN(_07391_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][14] ), .QN(_07392_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][13] ), .QN(_07393_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][12] ), .QN(_07394_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][29] ), .QN(_07395_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][11] ), .QN(_07396_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][10] ), .QN(_07397_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][9] ), .QN(_07398_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][8] ), .QN(_07399_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][7] ), .QN(_07400_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][6] ), .QN(_07401_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][5] ), .QN(_07402_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][4] ), .QN(_07403_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][3] ), .QN(_07404_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][2] ), .QN(_07405_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][28] ), .QN(_07406_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][1] ), .QN(_07407_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][0] ), .QN(_07408_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][27] ), .QN(_07409_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][26] ), .QN(_07410_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][25] ), .QN(_07411_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][24] ), .QN(_07412_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][23] ), .QN(_07413_ ) );
DFF_X1 \u_icache.cblocks[2]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06652_ ), .Q(\u_icache.cblocks[2][22] ), .QN(_07414_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][31] ), .QN(_07415_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][30] ), .QN(_07416_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][21] ), .QN(_07417_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][20] ), .QN(_07418_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][19] ), .QN(_07419_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][18] ), .QN(_07420_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][17] ), .QN(_07421_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][16] ), .QN(_07422_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][15] ), .QN(_07423_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][14] ), .QN(_07424_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][13] ), .QN(_07425_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][12] ), .QN(_07426_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][29] ), .QN(_07427_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][11] ), .QN(_07428_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][10] ), .QN(_07429_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][9] ), .QN(_07430_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][8] ), .QN(_07431_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][7] ), .QN(_07432_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][6] ), .QN(_07433_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][5] ), .QN(_07434_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][4] ), .QN(_07435_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][3] ), .QN(_07436_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][2] ), .QN(_07437_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][28] ), .QN(_07438_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][1] ), .QN(_07439_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][0] ), .QN(_07440_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][27] ), .QN(_07441_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][26] ), .QN(_07442_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][25] ), .QN(_07443_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][24] ), .QN(_07444_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][23] ), .QN(_07445_ ) );
DFF_X1 \u_icache.cblocks[3]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06651_ ), .Q(\u_icache.cblocks[3][22] ), .QN(_07446_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][31] ), .QN(_07447_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][30] ), .QN(_07448_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][21] ), .QN(_07449_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][20] ), .QN(_07450_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][19] ), .QN(_07451_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][18] ), .QN(_07452_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][17] ), .QN(_07453_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][16] ), .QN(_07454_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][15] ), .QN(_07455_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][14] ), .QN(_07456_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][13] ), .QN(_07457_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][12] ), .QN(_07458_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][29] ), .QN(_07459_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][11] ), .QN(_07460_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][10] ), .QN(_07461_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][9] ), .QN(_07462_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][8] ), .QN(_07463_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][7] ), .QN(_07464_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][6] ), .QN(_07465_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][5] ), .QN(_07466_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][4] ), .QN(_07467_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][3] ), .QN(_07468_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][2] ), .QN(_07469_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][28] ), .QN(_07470_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][1] ), .QN(_07471_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][0] ), .QN(_07472_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][27] ), .QN(_07473_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][26] ), .QN(_07474_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][25] ), .QN(_07475_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][24] ), .QN(_07476_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][23] ), .QN(_07477_ ) );
DFF_X1 \u_icache.cblocks[4]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06650_ ), .Q(\u_icache.cblocks[4][22] ), .QN(_07478_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][31] ), .QN(_07479_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][30] ), .QN(_07480_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][21] ), .QN(_07481_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][20] ), .QN(_07482_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][19] ), .QN(_07483_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][18] ), .QN(_07484_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][17] ), .QN(_07485_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][16] ), .QN(_07486_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][15] ), .QN(_07487_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][14] ), .QN(_07488_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][13] ), .QN(_07489_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][12] ), .QN(_07490_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][29] ), .QN(_07491_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][11] ), .QN(_07492_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][10] ), .QN(_07493_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][9] ), .QN(_07494_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][8] ), .QN(_07495_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][7] ), .QN(_07496_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][6] ), .QN(_07497_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][5] ), .QN(_07498_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][4] ), .QN(_07499_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][3] ), .QN(_07500_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][2] ), .QN(_07501_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][28] ), .QN(_07502_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][1] ), .QN(_07503_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][0] ), .QN(_07504_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][27] ), .QN(_07505_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][26] ), .QN(_07506_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][25] ), .QN(_07507_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][24] ), .QN(_07508_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][23] ), .QN(_07509_ ) );
DFF_X1 \u_icache.cblocks[5]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06649_ ), .Q(\u_icache.cblocks[5][22] ), .QN(_07510_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][31] ), .QN(_07511_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][30] ), .QN(_07512_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][21] ), .QN(_07513_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][20] ), .QN(_07514_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][19] ), .QN(_07515_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][18] ), .QN(_07516_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][17] ), .QN(_07517_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][16] ), .QN(_07518_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][15] ), .QN(_07519_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][14] ), .QN(_07520_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][13] ), .QN(_07521_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][12] ), .QN(_07522_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][29] ), .QN(_07523_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][11] ), .QN(_07524_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][10] ), .QN(_07525_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][9] ), .QN(_07526_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][8] ), .QN(_07527_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][7] ), .QN(_07528_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][6] ), .QN(_07529_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][5] ), .QN(_07530_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][4] ), .QN(_07531_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][3] ), .QN(_07532_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][2] ), .QN(_07533_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][28] ), .QN(_07534_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][1] ), .QN(_07535_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][0] ), .QN(_07536_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][27] ), .QN(_07537_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][26] ), .QN(_07538_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][25] ), .QN(_07539_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][24] ), .QN(_07540_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][23] ), .QN(_07541_ ) );
DFF_X1 \u_icache.cblocks[6]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06648_ ), .Q(\u_icache.cblocks[6][22] ), .QN(_07542_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q ( .D(\ac_data [31] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][31] ), .QN(_07543_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_1 ( .D(\ac_data [30] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][30] ), .QN(_07544_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_10 ( .D(\ac_data [21] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][21] ), .QN(_07545_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_11 ( .D(\ac_data [20] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][20] ), .QN(_07546_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_12 ( .D(\ac_data [19] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][19] ), .QN(_07547_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_13 ( .D(\ac_data [18] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][18] ), .QN(_07548_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_14 ( .D(\ac_data [17] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][17] ), .QN(_07549_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_15 ( .D(\ac_data [16] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][16] ), .QN(_07550_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_16 ( .D(\ac_data [15] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][15] ), .QN(_07551_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_17 ( .D(\ac_data [14] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][14] ), .QN(_07552_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_18 ( .D(\ac_data [13] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][13] ), .QN(_07553_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_19 ( .D(\ac_data [12] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][12] ), .QN(_07554_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_2 ( .D(\ac_data [29] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][29] ), .QN(_07555_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_20 ( .D(\ac_data [11] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][11] ), .QN(_07556_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_21 ( .D(\ac_data [10] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][10] ), .QN(_07557_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_22 ( .D(\ac_data [9] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][9] ), .QN(_07558_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_23 ( .D(\ac_data [8] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][8] ), .QN(_07559_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_24 ( .D(\ac_data [7] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][7] ), .QN(_07560_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_25 ( .D(\ac_data [6] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][6] ), .QN(_07561_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_26 ( .D(\ac_data [5] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][5] ), .QN(_07562_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_27 ( .D(\ac_data [4] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][4] ), .QN(_07563_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_28 ( .D(\ac_data [3] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][3] ), .QN(_07564_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_29 ( .D(\ac_data [2] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][2] ), .QN(_07565_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_3 ( .D(\ac_data [28] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][28] ), .QN(_07566_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_30 ( .D(\ac_data [1] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][1] ), .QN(_07567_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_31 ( .D(\ac_data [0] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][0] ), .QN(_07568_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_4 ( .D(\ac_data [27] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][27] ), .QN(_07569_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_5 ( .D(\ac_data [26] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][26] ), .QN(_07570_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_6 ( .D(\ac_data [25] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][25] ), .QN(_07571_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_7 ( .D(\ac_data [24] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][24] ), .QN(_07572_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_8 ( .D(\ac_data [23] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][23] ), .QN(_07573_ ) );
DFF_X1 \u_icache.cblocks[7]_$_DFFE_PP__Q_9 ( .D(\ac_data [22] ), .CK(_06647_ ), .Q(\u_icache.cblocks[7][22] ), .QN(_06873_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q ( .D(_00382_ ), .CK(_06646_ ), .Q(\cf_inst [31] ), .QN(_06872_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_1 ( .D(_00383_ ), .CK(_06646_ ), .Q(\cf_inst [30] ), .QN(_06871_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_10 ( .D(_00384_ ), .CK(_06646_ ), .Q(\cf_inst [21] ), .QN(_06870_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_11 ( .D(_00385_ ), .CK(_06646_ ), .Q(\cf_inst [20] ), .QN(_06869_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_12 ( .D(_00386_ ), .CK(_06646_ ), .Q(\cf_inst [19] ), .QN(_06868_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_13 ( .D(_00387_ ), .CK(_06646_ ), .Q(\cf_inst [18] ), .QN(_06867_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_14 ( .D(_00388_ ), .CK(_06646_ ), .Q(\cf_inst [17] ), .QN(_06866_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_15 ( .D(_00389_ ), .CK(_06646_ ), .Q(\cf_inst [16] ), .QN(_06865_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_16 ( .D(_00390_ ), .CK(_06646_ ), .Q(\cf_inst [15] ), .QN(_06864_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_17 ( .D(_00391_ ), .CK(_06646_ ), .Q(\cf_inst [14] ), .QN(_06863_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_18 ( .D(_00392_ ), .CK(_06646_ ), .Q(\cf_inst [13] ), .QN(_06862_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_19 ( .D(_00393_ ), .CK(_06646_ ), .Q(\cf_inst [12] ), .QN(_06861_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_2 ( .D(_00394_ ), .CK(_06646_ ), .Q(\cf_inst [29] ), .QN(_06860_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_20 ( .D(_00395_ ), .CK(_06646_ ), .Q(\cf_inst [11] ), .QN(_06859_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_21 ( .D(_00396_ ), .CK(_06646_ ), .Q(\cf_inst [10] ), .QN(_06858_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_22 ( .D(_00397_ ), .CK(_06646_ ), .Q(\cf_inst [9] ), .QN(_06857_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_23 ( .D(_00398_ ), .CK(_06646_ ), .Q(\cf_inst [8] ), .QN(_06856_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_24 ( .D(_00399_ ), .CK(_06646_ ), .Q(\cf_inst [7] ), .QN(_06855_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_25 ( .D(_00400_ ), .CK(_06646_ ), .Q(\cf_inst [6] ), .QN(_06854_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_26 ( .D(_00401_ ), .CK(_06646_ ), .Q(\cf_inst [5] ), .QN(_06853_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_27 ( .D(_00402_ ), .CK(_06646_ ), .Q(\cf_inst [4] ), .QN(_06852_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_28 ( .D(_00403_ ), .CK(_06646_ ), .Q(\cf_inst [3] ), .QN(_06851_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_29 ( .D(_00404_ ), .CK(_06646_ ), .Q(\cf_inst [2] ), .QN(_06850_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_3 ( .D(_00405_ ), .CK(_06646_ ), .Q(\cf_inst [28] ), .QN(_06849_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_30 ( .D(_00406_ ), .CK(_06646_ ), .Q(\cf_inst [1] ), .QN(_06848_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_31 ( .D(_00407_ ), .CK(_06646_ ), .Q(\cf_inst [0] ), .QN(_06847_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_4 ( .D(_00408_ ), .CK(_06646_ ), .Q(\cf_inst [27] ), .QN(_06846_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_5 ( .D(_00409_ ), .CK(_06646_ ), .Q(\cf_inst [26] ), .QN(_06845_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_6 ( .D(_00410_ ), .CK(_06646_ ), .Q(\cf_inst [25] ), .QN(_06844_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_7 ( .D(_00411_ ), .CK(_06646_ ), .Q(\cf_inst [24] ), .QN(_06843_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_8 ( .D(_00412_ ), .CK(_06646_ ), .Q(\cf_inst [23] ), .QN(_06842_ ) );
DFF_X1 \u_icache.cdata_$_SDFFE_PP0P__Q_9 ( .D(_00413_ ), .CK(_06646_ ), .Q(\cf_inst [22] ), .QN(_06841_ ) );
DFF_X1 \u_icache.chvalid_$_SDFFE_PP0P__Q ( .D(_00414_ ), .CK(_06645_ ), .Q(icah_valid ), .QN(\u_lsu.reading_$_NOR__B_A_$_MUX__Y_B ) );
DFF_X1 \u_icache.count_$_SDFFE_PP0P__Q ( .D(_00415_ ), .CK(_06644_ ), .Q(\u_icache.count [2] ), .QN(_06840_ ) );
DFF_X1 \u_icache.count_$_SDFFE_PP0P__Q_1 ( .D(_00416_ ), .CK(_06644_ ), .Q(\u_icache.count [1] ), .QN(_06839_ ) );
DFF_X1 \u_icache.count_$_SDFFE_PP0P__Q_2 ( .D(_00417_ ), .CK(_06644_ ), .Q(\u_icache.count [0] ), .QN(\u_icache.count_$_NOT__A_Y ) );
DFF_X1 \u_icache.cready_$_SDFF_PP0__Q ( .D(_00418_ ), .CK(clock ), .Q(ifu_ready ), .QN(_07574_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q ( .D(\fc_addr [31] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][26] ), .QN(_06838_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_1 ( .D(\fc_addr [30] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][25] ), .QN(_07575_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_10 ( .D(\fc_addr [21] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][16] ), .QN(_07576_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_11 ( .D(\fc_addr [20] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][15] ), .QN(_07577_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_12 ( .D(\fc_addr [19] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][14] ), .QN(_07578_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_13 ( .D(\fc_addr [18] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][13] ), .QN(_07579_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_14 ( .D(\fc_addr [17] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][12] ), .QN(_07580_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_15 ( .D(\fc_addr [16] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][11] ), .QN(_07581_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_16 ( .D(\fc_addr [15] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][10] ), .QN(_07582_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_17 ( .D(\fc_addr [14] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][9] ), .QN(_07583_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_18 ( .D(\fc_addr [13] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][8] ), .QN(_07584_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_19 ( .D(\fc_addr [12] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][7] ), .QN(_07585_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_2 ( .D(\fc_addr [29] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][24] ), .QN(_07586_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_20 ( .D(\fc_addr [11] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][6] ), .QN(_07587_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_21 ( .D(\fc_addr [10] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][5] ), .QN(_07588_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_22 ( .D(\fc_addr [9] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][4] ), .QN(_07589_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_23 ( .D(\fc_addr [8] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][3] ), .QN(_07590_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_24 ( .D(\fc_addr [7] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][2] ), .QN(_07591_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_25 ( .D(\fc_addr [6] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][1] ), .QN(_07592_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_26 ( .D(\fc_addr [5] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][0] ), .QN(_07593_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_3 ( .D(\fc_addr [28] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][23] ), .QN(_07594_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_4 ( .D(\fc_addr [27] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][22] ), .QN(_07595_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_5 ( .D(\fc_addr [26] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][21] ), .QN(_07596_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_6 ( .D(\fc_addr [25] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][20] ), .QN(_07597_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_7 ( .D(\fc_addr [24] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][19] ), .QN(_07598_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_8 ( .D(\fc_addr [23] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][18] ), .QN(_07599_ ) );
DFF_X1 \u_icache.ctags[0]_$_DFFE_PP__Q_9 ( .D(\fc_addr [22] ), .CK(_06643_ ), .Q(\u_icache.ctags[0][17] ), .QN(_07600_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q ( .D(\fc_addr [31] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][26] ), .QN(_07601_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_1 ( .D(\fc_addr [30] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][25] ), .QN(_07602_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_10 ( .D(\fc_addr [21] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][16] ), .QN(_07603_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_11 ( .D(\fc_addr [20] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][15] ), .QN(_07604_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_12 ( .D(\fc_addr [19] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][14] ), .QN(_07605_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_13 ( .D(\fc_addr [18] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][13] ), .QN(_07606_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_14 ( .D(\fc_addr [17] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][12] ), .QN(_07607_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_15 ( .D(\fc_addr [16] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][11] ), .QN(_07608_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_16 ( .D(\fc_addr [15] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][10] ), .QN(_07609_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_17 ( .D(\fc_addr [14] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][9] ), .QN(_07610_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_18 ( .D(\fc_addr [13] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][8] ), .QN(_07611_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_19 ( .D(\fc_addr [12] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][7] ), .QN(_07612_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_2 ( .D(\fc_addr [29] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][24] ), .QN(_07613_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_20 ( .D(\fc_addr [11] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][6] ), .QN(_07614_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_21 ( .D(\fc_addr [10] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][5] ), .QN(_07615_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_22 ( .D(\fc_addr [9] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][4] ), .QN(_07616_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_23 ( .D(\fc_addr [8] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][3] ), .QN(_07617_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_24 ( .D(\fc_addr [7] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][2] ), .QN(_07618_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_25 ( .D(\fc_addr [6] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][1] ), .QN(_07619_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_26 ( .D(\fc_addr [5] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][0] ), .QN(_07620_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_3 ( .D(\fc_addr [28] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][23] ), .QN(_07621_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_4 ( .D(\fc_addr [27] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][22] ), .QN(_07622_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_5 ( .D(\fc_addr [26] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][21] ), .QN(_07623_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_6 ( .D(\fc_addr [25] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][20] ), .QN(_07624_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_7 ( .D(\fc_addr [24] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][19] ), .QN(_07625_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_8 ( .D(\fc_addr [23] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][18] ), .QN(_07626_ ) );
DFF_X1 \u_icache.ctags[1]_$_DFFE_PP__Q_9 ( .D(\fc_addr [22] ), .CK(_06642_ ), .Q(\u_icache.ctags[1][17] ), .QN(_06837_ ) );
DFF_X1 \u_icache.cvalids_$_SDFFE_PP0P__Q ( .D(_00419_ ), .CK(_06641_ ), .Q(\u_icache.cvalids [1] ), .QN(_06836_ ) );
DFF_X1 \u_icache.cvalids_$_SDFFE_PP0P__Q_1 ( .D(_00420_ ), .CK(_06641_ ), .Q(\u_icache.cvalids [0] ), .QN(_06835_ ) );
DFF_X1 \u_icache.ended_$_SDFFE_PP0P__Q ( .D(_00421_ ), .CK(_06640_ ), .Q(\u_icache.ended ), .QN(_06834_ ) );
DFF_X1 \u_idu.decode_ok_$_SDFFE_PP0P__Q ( .D(_00422_ ), .CK(_06639_ ), .Q(exe_valid ), .QN(_06833_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q ( .D(_00423_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [31] ), .QN(_06832_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_1 ( .D(_00424_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [30] ), .QN(\u_exu.opt_$_NOR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_10 ( .D(_00425_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [21] ), .QN(_06831_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_11 ( .D(_00426_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [20] ), .QN(\u_idu.errmux_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_NAND__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_12 ( .D(_00427_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [19] ), .QN(_06830_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_13 ( .D(_00428_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [18] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_14 ( .D(_00429_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [17] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_1_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_15 ( .D(_00430_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [16] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_2_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_16 ( .D(_00431_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [15] ), .QN(_06829_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_17 ( .D(_00432_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [14] ), .QN(de_ard_$_NOR__Y_1_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_18 ( .D(_00433_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [13] ), .QN(de_ard_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_19 ( .D(_00434_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [12] ), .QN(\u_exu.alu_ctrl_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_2 ( .D(_00435_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [29] ), .QN(_06828_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_20 ( .D(_00436_ ), .CK(_06638_ ), .Q(\u_idu.imm_branch [4] ), .QN(_06827_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_21 ( .D(_00437_ ), .CK(_06638_ ), .Q(\u_idu.imm_branch [3] ), .QN(_06826_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_22 ( .D(_00438_ ), .CK(_06638_ ), .Q(\u_idu.imm_branch [2] ), .QN(_06825_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_23 ( .D(_00439_ ), .CK(_06638_ ), .Q(\u_idu.imm_branch [1] ), .QN(_06824_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_24 ( .D(_00440_ ), .CK(_06638_ ), .Q(\u_idu.imm_branch [11] ), .QN(_06823_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_25 ( .D(_00441_ ), .CK(_06638_ ), .Q(\u_idu.inst [6] ), .QN(\u_exu.opt_$_NOR__Y_2_A_$_ANDNOT__Y_A_$_ANDNOT__A_B_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_A_$_OR__A_B ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_26 ( .D(_00442_ ), .CK(_06638_ ), .Q(\u_idu.inst [5] ), .QN(_06822_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_27 ( .D(_00443_ ), .CK(_06638_ ), .Q(\u_idu.inst [4] ), .QN(_06821_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_28 ( .D(_00444_ ), .CK(_06638_ ), .Q(\u_idu.inst [3] ), .QN(_06820_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_29 ( .D(_00445_ ), .CK(_06638_ ), .Q(\u_idu.inst [2] ), .QN(_06819_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_3 ( .D(_00446_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [28] ), .QN(_06818_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_30 ( .D(_00447_ ), .CK(_06638_ ), .Q(\u_idu.inst [1] ), .QN(_06817_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_31 ( .D(_00448_ ), .CK(_06638_ ), .Q(\u_idu.inst [0] ), .QN(_06816_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_4 ( .D(_00449_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [27] ), .QN(_06815_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_5 ( .D(_00450_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [26] ), .QN(_06814_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_6 ( .D(_00451_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [25] ), .QN(_06813_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_7 ( .D(_00452_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [24] ), .QN(_06812_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_8 ( .D(_00453_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [23] ), .QN(_06811_ ) );
DFF_X1 \u_idu.inst_$_SDFFE_PP0P__Q_9 ( .D(_00454_ ), .CK(_06638_ ), .Q(\u_idu.imm_auipc_lui [22] ), .QN(_06810_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q ( .D(_00455_ ), .CK(_06638_ ), .Q(\de_pc [31] ), .QN(_06809_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00456_ ), .CK(_06638_ ), .Q(\de_pc [30] ), .QN(_06808_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00457_ ), .CK(_06638_ ), .Q(\de_pc [21] ), .QN(_06807_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00458_ ), .CK(_06638_ ), .Q(\de_pc [20] ), .QN(_06806_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00459_ ), .CK(_06638_ ), .Q(\de_pc [19] ), .QN(_06805_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00460_ ), .CK(_06638_ ), .Q(\de_pc [18] ), .QN(_06804_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00461_ ), .CK(_06638_ ), .Q(\de_pc [17] ), .QN(_06803_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00462_ ), .CK(_06638_ ), .Q(\de_pc [16] ), .QN(_06802_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00463_ ), .CK(_06638_ ), .Q(\de_pc [15] ), .QN(_06801_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00464_ ), .CK(_06638_ ), .Q(\de_pc [14] ), .QN(_06800_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00465_ ), .CK(_06638_ ), .Q(\de_pc [13] ), .QN(_06799_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00466_ ), .CK(_06638_ ), .Q(\de_pc [12] ), .QN(_06798_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00467_ ), .CK(_06638_ ), .Q(\de_pc [29] ), .QN(_06797_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00468_ ), .CK(_06638_ ), .Q(\de_pc [11] ), .QN(_06796_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00469_ ), .CK(_06638_ ), .Q(\de_pc [10] ), .QN(_06795_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00470_ ), .CK(_06638_ ), .Q(\de_pc [9] ), .QN(_06794_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00471_ ), .CK(_06638_ ), .Q(\de_pc [8] ), .QN(_06793_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00472_ ), .CK(_06638_ ), .Q(\de_pc [7] ), .QN(_06792_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00473_ ), .CK(_06638_ ), .Q(\de_pc [6] ), .QN(_06791_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00474_ ), .CK(_06638_ ), .Q(\de_pc [5] ), .QN(_06790_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00475_ ), .CK(_06638_ ), .Q(\de_pc [4] ), .QN(_06789_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00476_ ), .CK(_06638_ ), .Q(\de_pc [3] ), .QN(_06788_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00477_ ), .CK(_06638_ ), .Q(\de_pc [2] ), .QN(_06787_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00478_ ), .CK(_06638_ ), .Q(\de_pc [28] ), .QN(_06786_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00479_ ), .CK(_06638_ ), .Q(\de_pc [1] ), .QN(_06785_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_31 ( .D(_00480_ ), .CK(_06638_ ), .Q(\de_pc [0] ), .QN(_06784_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00481_ ), .CK(_06638_ ), .Q(\de_pc [27] ), .QN(_06783_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00482_ ), .CK(_06638_ ), .Q(\de_pc [26] ), .QN(_06782_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00483_ ), .CK(_06638_ ), .Q(\de_pc [25] ), .QN(_06781_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00484_ ), .CK(_06638_ ), .Q(\de_pc [24] ), .QN(_06780_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00485_ ), .CK(_06638_ ), .Q(\de_pc [23] ), .QN(_06779_ ) );
DFF_X1 \u_idu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00486_ ), .CK(_06638_ ), .Q(\de_pc [22] ), .QN(_06778_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q ( .D(_00487_ ), .CK(_06637_ ), .Q(\fd_inst [31] ), .QN(_06777_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_1 ( .D(_00488_ ), .CK(_06637_ ), .Q(\fd_inst [30] ), .QN(_06776_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_10 ( .D(_00489_ ), .CK(_06637_ ), .Q(\fd_inst [21] ), .QN(_06775_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_11 ( .D(_00490_ ), .CK(_06637_ ), .Q(\fd_inst [20] ), .QN(_06774_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_12 ( .D(_00491_ ), .CK(_06637_ ), .Q(\fd_inst [19] ), .QN(_06773_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_13 ( .D(_00492_ ), .CK(_06637_ ), .Q(\fd_inst [18] ), .QN(_06772_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_14 ( .D(_00493_ ), .CK(_06637_ ), .Q(\fd_inst [17] ), .QN(_06771_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_15 ( .D(_00494_ ), .CK(_06637_ ), .Q(\fd_inst [16] ), .QN(_06770_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_16 ( .D(_00495_ ), .CK(_06637_ ), .Q(\fd_inst [15] ), .QN(_06769_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_17 ( .D(_00496_ ), .CK(_06637_ ), .Q(\fd_inst [14] ), .QN(_06768_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_18 ( .D(_00497_ ), .CK(_06637_ ), .Q(\fd_inst [13] ), .QN(_06767_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_19 ( .D(_00498_ ), .CK(_06637_ ), .Q(\fd_inst [12] ), .QN(_06766_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_2 ( .D(_00499_ ), .CK(_06637_ ), .Q(\fd_inst [29] ), .QN(_06765_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_20 ( .D(_00500_ ), .CK(_06637_ ), .Q(\fd_inst [11] ), .QN(_06764_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_21 ( .D(_00501_ ), .CK(_06637_ ), .Q(\fd_inst [10] ), .QN(_06763_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_22 ( .D(_00502_ ), .CK(_06637_ ), .Q(\fd_inst [9] ), .QN(_06762_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_23 ( .D(_00503_ ), .CK(_06637_ ), .Q(\fd_inst [8] ), .QN(_06761_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_24 ( .D(_00504_ ), .CK(_06637_ ), .Q(\fd_inst [7] ), .QN(_06760_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_25 ( .D(_00505_ ), .CK(_06637_ ), .Q(\fd_inst [6] ), .QN(_06759_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_26 ( .D(_00506_ ), .CK(_06637_ ), .Q(\fd_inst [5] ), .QN(_06758_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_27 ( .D(_00507_ ), .CK(_06637_ ), .Q(\fd_inst [4] ), .QN(_06757_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_28 ( .D(_00508_ ), .CK(_06637_ ), .Q(\fd_inst [3] ), .QN(_06756_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_29 ( .D(_00509_ ), .CK(_06637_ ), .Q(\fd_inst [2] ), .QN(_06755_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_3 ( .D(_00510_ ), .CK(_06637_ ), .Q(\fd_inst [28] ), .QN(_06754_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_30 ( .D(_00511_ ), .CK(_06637_ ), .Q(\fd_inst [1] ), .QN(_06753_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_31 ( .D(_00512_ ), .CK(_06637_ ), .Q(\fd_inst [0] ), .QN(_06752_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_4 ( .D(_00513_ ), .CK(_06637_ ), .Q(\fd_inst [27] ), .QN(_06751_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_5 ( .D(_00514_ ), .CK(_06637_ ), .Q(\fd_inst [26] ), .QN(_06750_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_6 ( .D(_00515_ ), .CK(_06637_ ), .Q(\fd_inst [25] ), .QN(_06749_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_7 ( .D(_00516_ ), .CK(_06637_ ), .Q(\fd_inst [24] ), .QN(_06748_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_8 ( .D(_00517_ ), .CK(_06637_ ), .Q(\fd_inst [23] ), .QN(_06747_ ) );
DFF_X1 \u_ifu.inst_$_SDFFE_PP0P__Q_9 ( .D(_00518_ ), .CK(_06637_ ), .Q(\fd_inst [22] ), .QN(_06746_ ) );
DFF_X1 \u_ifu.inst_ok_$_SDFFE_PP0P__Q ( .D(_00519_ ), .CK(_06636_ ), .Q(idu_ready ), .QN(_06745_ ) );
DFF_X1 \u_ifu.jpc_ok_$_SDFFE_PP0P__Q ( .D(_00520_ ), .CK(_06635_ ), .Q(\u_ifu.jpc_ok ), .QN(\u_ifu.jpc_ok_$_NOT__A_Y ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q ( .D(_00521_ ), .CK(_06634_ ), .Q(\fc_addr [30] ), .QN(_06744_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_1 ( .D(_00522_ ), .CK(_06634_ ), .Q(\fc_addr [29] ), .QN(_06743_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_10 ( .D(_00523_ ), .CK(_06634_ ), .Q(\fc_addr [20] ), .QN(_06742_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_11 ( .D(_00524_ ), .CK(_06634_ ), .Q(\fc_addr [19] ), .QN(_06741_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_12 ( .D(_00525_ ), .CK(_06634_ ), .Q(\fc_addr [18] ), .QN(_06740_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_13 ( .D(_00526_ ), .CK(_06634_ ), .Q(\fc_addr [17] ), .QN(_06739_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_14 ( .D(_00527_ ), .CK(_06634_ ), .Q(\fc_addr [16] ), .QN(_06738_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_15 ( .D(_00528_ ), .CK(_06634_ ), .Q(\fc_addr [15] ), .QN(_06737_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_16 ( .D(_00529_ ), .CK(_06634_ ), .Q(\fc_addr [14] ), .QN(_06736_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_17 ( .D(_00530_ ), .CK(_06634_ ), .Q(\fc_addr [13] ), .QN(_06735_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_18 ( .D(_00531_ ), .CK(_06634_ ), .Q(\fc_addr [12] ), .QN(_06734_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_19 ( .D(_00532_ ), .CK(_06634_ ), .Q(\fc_addr [11] ), .QN(_06733_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_2 ( .D(_00533_ ), .CK(_06634_ ), .Q(\fc_addr [28] ), .QN(_06732_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_20 ( .D(_00534_ ), .CK(_06634_ ), .Q(\fc_addr [10] ), .QN(_06731_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_21 ( .D(_00535_ ), .CK(_06634_ ), .Q(\fc_addr [9] ), .QN(_06730_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_22 ( .D(_00536_ ), .CK(_06634_ ), .Q(\fc_addr [8] ), .QN(_06729_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_23 ( .D(_00537_ ), .CK(_06634_ ), .Q(\fc_addr [7] ), .QN(_06728_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_24 ( .D(_00538_ ), .CK(_06634_ ), .Q(\fc_addr [6] ), .QN(_06727_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_25 ( .D(_00539_ ), .CK(_06634_ ), .Q(\fc_addr [5] ), .QN(_06726_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_26 ( .D(_00540_ ), .CK(_06634_ ), .Q(\fc_addr [4] ), .QN(\u_ifu.pc_$_SDFFE_PP0N__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D ( .D(_00542_ ), .CK(clock ), .Q(\u_ifu.pc_$_SDFFE_PP0N__Q_26_D_$_MUX__A_Y_$_SDFF_PP0__D_Q ), .QN(_06724_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_27 ( .D(_00541_ ), .CK(_06634_ ), .Q(\fc_addr [3] ), .QN(_06725_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_28 ( .D(_00543_ ), .CK(_06634_ ), .Q(\fc_addr [2] ), .QN(\u_ifu.pc_$_SDFFE_PP0N__Q_28_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_3 ( .D(_00544_ ), .CK(_06634_ ), .Q(\fc_addr [27] ), .QN(_06723_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_4 ( .D(_00545_ ), .CK(_06634_ ), .Q(\fc_addr [26] ), .QN(_06722_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_5 ( .D(_00546_ ), .CK(_06634_ ), .Q(\fc_addr [25] ), .QN(_06721_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_6 ( .D(_00547_ ), .CK(_06634_ ), .Q(\fc_addr [24] ), .QN(_06720_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_7 ( .D(_00548_ ), .CK(_06634_ ), .Q(\fc_addr [23] ), .QN(_06719_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_8 ( .D(_00549_ ), .CK(_06634_ ), .Q(\fc_addr [22] ), .QN(_06718_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0N__Q_9 ( .D(_00550_ ), .CK(_06634_ ), .Q(\fc_addr [21] ), .QN(_06717_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0P__Q ( .D(_00551_ ), .CK(_06633_ ), .Q(\fc_addr [1] ), .QN(_06716_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00552_ ), .CK(_06633_ ), .Q(\fc_addr [0] ), .QN(_06715_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP1N__Q ( .D(_00553_ ), .CK(_06634_ ), .Q(\fc_addr [31] ), .QN(_06714_ ) );
DFF_X1 \u_lsu.arvalid_$_SDFFE_PP0P__Q ( .D(_00554_ ), .CK(_06632_ ), .Q(\u_lsu.arvalid ), .QN(_06713_ ) );
DFF_X1 \u_lsu.awvalid_$_SDFFE_PP0P__Q ( .D(_00555_ ), .CK(_06631_ ), .Q(io_master_awvalid ), .QN(_06712_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q ( .D(_00556_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [7] ), .QN(_06711_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_1 ( .D(_00557_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [6] ), .QN(_06710_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_2 ( .D(_00558_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [5] ), .QN(_06709_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_3 ( .D(_00559_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [4] ), .QN(_06708_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_4 ( .D(_00560_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [3] ), .QN(_06707_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_5 ( .D(_00561_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [2] ), .QN(_06706_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_6 ( .D(_00562_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [1] ), .QN(_06705_ ) );
DFF_X1 \u_lsu.rcount_$_SDFFE_PP0P__Q_7 ( .D(_00563_ ), .CK(_06630_ ), .Q(\u_lsu.rcount [0] ), .QN(_06704_ ) );
DFF_X1 \u_lsu.reading_$_SDFFE_PP0P__Q ( .D(_00554_ ), .CK(_06629_ ), .Q(\u_lsu.reading ), .QN(_06703_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q ( .D(_00564_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [63] ), .QN(_06701_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_1 ( .D(_00565_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [62] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_10 ( .D(_00566_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [53] ), .QN(_06700_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_11 ( .D(_00567_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [52] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_10_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_12 ( .D(_00568_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [51] ), .QN(_06699_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_13 ( .D(_00569_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [50] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_12_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_14 ( .D(_00570_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [49] ), .QN(_06698_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_15 ( .D(_00571_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [48] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_14_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_16 ( .D(_00572_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [47] ), .QN(_06697_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_17 ( .D(_00573_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [46] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_16_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_18 ( .D(_00574_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [45] ), .QN(_06696_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_19 ( .D(_00575_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [44] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_18_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_2 ( .D(_00576_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [61] ), .QN(_06695_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_20 ( .D(_00577_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [43] ), .QN(_06694_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_21 ( .D(_00578_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [42] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_20_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_22 ( .D(_00579_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [41] ), .QN(_06693_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_23 ( .D(_00580_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [40] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_22_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_24 ( .D(_00581_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [39] ), .QN(_06692_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_25 ( .D(_00582_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [38] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_24_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_26 ( .D(_00583_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [37] ), .QN(_06691_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_27 ( .D(_00584_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [36] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_26_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_28 ( .D(_00585_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [35] ), .QN(_06690_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_29 ( .D(_00586_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [34] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_28_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_3 ( .D(_00587_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [60] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_2_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_30 ( .D(_00588_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [33] ), .QN(_06689_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_31 ( .D(_00589_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [32] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_32 ( .D(_00590_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [31] ), .QN(_06688_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_33 ( .D(_00591_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [30] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_31_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_34 ( .D(_00592_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [29] ), .QN(_06687_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_35 ( .D(_00593_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [28] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_33_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_36 ( .D(_00594_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [27] ), .QN(_06686_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_37 ( .D(_00595_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [26] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_35_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_38 ( .D(_00596_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [25] ), .QN(_06685_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_39 ( .D(_00597_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [24] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_37_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_4 ( .D(_00598_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [59] ), .QN(_06684_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_40 ( .D(_00599_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [23] ), .QN(_06683_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_41 ( .D(_00600_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [22] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_39_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_42 ( .D(_00601_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [21] ), .QN(_06682_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_43 ( .D(_00602_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [20] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_41_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_44 ( .D(_00603_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [19] ), .QN(_06681_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_45 ( .D(_00604_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [18] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_43_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_46 ( .D(_00605_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [17] ), .QN(_06680_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_47 ( .D(_00606_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [16] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_45_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_48 ( .D(_00607_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [15] ), .QN(_06679_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_49 ( .D(_00608_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [14] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_47_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_5 ( .D(_00609_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [58] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_4_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_50 ( .D(_00610_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [13] ), .QN(_06678_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_51 ( .D(_00611_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [12] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_49_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_52 ( .D(_00612_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [11] ), .QN(_06677_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_53 ( .D(_00613_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [10] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_51_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_54 ( .D(_00614_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [9] ), .QN(_06676_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_55 ( .D(_00615_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [8] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_53_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_56 ( .D(_00616_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [7] ), .QN(_06675_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_57 ( .D(_00617_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [6] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_55_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_58 ( .D(_00618_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [5] ), .QN(_06674_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_59 ( .D(_00619_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [4] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_57_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_6 ( .D(_00620_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [57] ), .QN(_06673_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_60 ( .D(_00621_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [3] ), .QN(_06672_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_61 ( .D(_00622_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [2] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_59_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_62 ( .D(_00623_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [1] ), .QN(_06671_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63 ( .D(_00624_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [0] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_7 ( .D(_00625_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [56] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_6_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_8 ( .D(_00626_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [55] ), .QN(_06670_ ) );
DFF_X1 \u_lsu.u_clint.mtime_$_SDFF_PP0__Q_9 ( .D(_00627_ ), .CK(clock ), .Q(\u_lsu.u_clint.mtime [54] ), .QN(\u_lsu.u_clint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__B_A_$_ANDNOT__B_Y_$_XOR__A_Y_$_XOR__Y_8_A_$_ANDNOT__Y_B ) );
DFF_X1 \u_lsu.u_clint.tvalid_$_SDFF_PP0__Q ( .D(_00628_ ), .CK(clock ), .Q(\u_lsu.rvalid_clint ), .QN(\u_icache.chdata_$_ANDNOT__Y_23_B_$_OR__Y_A_$_AND__Y_B_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \u_lsu.wlast_$_SDFFE_PP0P__Q ( .D(_00555_ ), .CK(_06628_ ), .Q(io_master_wlast ), .QN(_06702_ ) );
DFF_X1 \u_lsu.writing_$_SDFFE_PP0P__Q ( .D(_00555_ ), .CK(_06627_ ), .Q(\u_lsu.writing ), .QN(_07627_ ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06626_ ), .Q(\u_reg.rf[10][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06626_ ), .Q(\u_reg.rf[10][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06626_ ), .Q(\u_reg.rf[10][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06626_ ), .Q(\u_reg.rf[10][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06626_ ), .Q(\u_reg.rf[10][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06626_ ), .Q(\u_reg.rf[10][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06626_ ), .Q(\u_reg.rf[10][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06626_ ), .Q(\u_reg.rf[10][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06626_ ), .Q(\u_reg.rf[10][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06626_ ), .Q(\u_reg.rf[10][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06626_ ), .Q(\u_reg.rf[10][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06626_ ), .Q(\u_reg.rf[10][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06626_ ), .Q(\u_reg.rf[10][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06626_ ), .Q(\u_reg.rf[10][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06626_ ), .Q(\u_reg.rf[10][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06626_ ), .Q(\u_reg.rf[10][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06626_ ), .Q(\u_reg.rf[10][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06626_ ), .Q(\u_reg.rf[10][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06626_ ), .Q(\u_reg.rf[10][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06626_ ), .Q(\u_reg.rf[10][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06626_ ), .Q(\u_reg.rf[10][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06626_ ), .Q(\u_reg.rf[10][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06626_ ), .Q(\u_reg.rf[10][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06626_ ), .Q(\u_reg.rf[10][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06626_ ), .Q(\u_reg.rf[10][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06626_ ), .Q(\u_reg.rf[10][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06626_ ), .Q(\u_reg.rf[10][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06626_ ), .Q(\u_reg.rf[10][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06626_ ), .Q(\u_reg.rf[10][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06626_ ), .Q(\u_reg.rf[10][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06626_ ), .Q(\u_reg.rf[10][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[10]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06626_ ), .Q(\u_reg.rf[10][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06625_ ), .Q(\u_reg.rf[11][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06625_ ), .Q(\u_reg.rf[11][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06625_ ), .Q(\u_reg.rf[11][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06625_ ), .Q(\u_reg.rf[11][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06625_ ), .Q(\u_reg.rf[11][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06625_ ), .Q(\u_reg.rf[11][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06625_ ), .Q(\u_reg.rf[11][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06625_ ), .Q(\u_reg.rf[11][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06625_ ), .Q(\u_reg.rf[11][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06625_ ), .Q(\u_reg.rf[11][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06625_ ), .Q(\u_reg.rf[11][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06625_ ), .Q(\u_reg.rf[11][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06625_ ), .Q(\u_reg.rf[11][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06625_ ), .Q(\u_reg.rf[11][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06625_ ), .Q(\u_reg.rf[11][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06625_ ), .Q(\u_reg.rf[11][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06625_ ), .Q(\u_reg.rf[11][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06625_ ), .Q(\u_reg.rf[11][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06625_ ), .Q(\u_reg.rf[11][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06625_ ), .Q(\u_reg.rf[11][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06625_ ), .Q(\u_reg.rf[11][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06625_ ), .Q(\u_reg.rf[11][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06625_ ), .Q(\u_reg.rf[11][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06625_ ), .Q(\u_reg.rf[11][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06625_ ), .Q(\u_reg.rf[11][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06625_ ), .Q(\u_reg.rf[11][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06625_ ), .Q(\u_reg.rf[11][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06625_ ), .Q(\u_reg.rf[11][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06625_ ), .Q(\u_reg.rf[11][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06625_ ), .Q(\u_reg.rf[11][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06625_ ), .Q(\u_reg.rf[11][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[11]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06625_ ), .Q(\u_reg.rf[11][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06624_ ), .Q(\u_reg.rf[12][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06624_ ), .Q(\u_reg.rf[12][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06624_ ), .Q(\u_reg.rf[12][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06624_ ), .Q(\u_reg.rf[12][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06624_ ), .Q(\u_reg.rf[12][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06624_ ), .Q(\u_reg.rf[12][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06624_ ), .Q(\u_reg.rf[12][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06624_ ), .Q(\u_reg.rf[12][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06624_ ), .Q(\u_reg.rf[12][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06624_ ), .Q(\u_reg.rf[12][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06624_ ), .Q(\u_reg.rf[12][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06624_ ), .Q(\u_reg.rf[12][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06624_ ), .Q(\u_reg.rf[12][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06624_ ), .Q(\u_reg.rf[12][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06624_ ), .Q(\u_reg.rf[12][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06624_ ), .Q(\u_reg.rf[12][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06624_ ), .Q(\u_reg.rf[12][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06624_ ), .Q(\u_reg.rf[12][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06624_ ), .Q(\u_reg.rf[12][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06624_ ), .Q(\u_reg.rf[12][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06624_ ), .Q(\u_reg.rf[12][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06624_ ), .Q(\u_reg.rf[12][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06624_ ), .Q(\u_reg.rf[12][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06624_ ), .Q(\u_reg.rf[12][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06624_ ), .Q(\u_reg.rf[12][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06624_ ), .Q(\u_reg.rf[12][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06624_ ), .Q(\u_reg.rf[12][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06624_ ), .Q(\u_reg.rf[12][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06624_ ), .Q(\u_reg.rf[12][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06624_ ), .Q(\u_reg.rf[12][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06624_ ), .Q(\u_reg.rf[12][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[12]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06624_ ), .Q(\u_reg.rf[12][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06623_ ), .Q(\u_reg.rf[13][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06623_ ), .Q(\u_reg.rf[13][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06623_ ), .Q(\u_reg.rf[13][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06623_ ), .Q(\u_reg.rf[13][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06623_ ), .Q(\u_reg.rf[13][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06623_ ), .Q(\u_reg.rf[13][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06623_ ), .Q(\u_reg.rf[13][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06623_ ), .Q(\u_reg.rf[13][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06623_ ), .Q(\u_reg.rf[13][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06623_ ), .Q(\u_reg.rf[13][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06623_ ), .Q(\u_reg.rf[13][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06623_ ), .Q(\u_reg.rf[13][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06623_ ), .Q(\u_reg.rf[13][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06623_ ), .Q(\u_reg.rf[13][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06623_ ), .Q(\u_reg.rf[13][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06623_ ), .Q(\u_reg.rf[13][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06623_ ), .Q(\u_reg.rf[13][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06623_ ), .Q(\u_reg.rf[13][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06623_ ), .Q(\u_reg.rf[13][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06623_ ), .Q(\u_reg.rf[13][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06623_ ), .Q(\u_reg.rf[13][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06623_ ), .Q(\u_reg.rf[13][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06623_ ), .Q(\u_reg.rf[13][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06623_ ), .Q(\u_reg.rf[13][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06623_ ), .Q(\u_reg.rf[13][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06623_ ), .Q(\u_reg.rf[13][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06623_ ), .Q(\u_reg.rf[13][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06623_ ), .Q(\u_reg.rf[13][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06623_ ), .Q(\u_reg.rf[13][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06623_ ), .Q(\u_reg.rf[13][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06623_ ), .Q(\u_reg.rf[13][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[13]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06623_ ), .Q(\u_reg.rf[13][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06622_ ), .Q(\u_reg.rf[14][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06622_ ), .Q(\u_reg.rf[14][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06622_ ), .Q(\u_reg.rf[14][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06622_ ), .Q(\u_reg.rf[14][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06622_ ), .Q(\u_reg.rf[14][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06622_ ), .Q(\u_reg.rf[14][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06622_ ), .Q(\u_reg.rf[14][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06622_ ), .Q(\u_reg.rf[14][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06622_ ), .Q(\u_reg.rf[14][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06622_ ), .Q(\u_reg.rf[14][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06622_ ), .Q(\u_reg.rf[14][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06622_ ), .Q(\u_reg.rf[14][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06622_ ), .Q(\u_reg.rf[14][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06622_ ), .Q(\u_reg.rf[14][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06622_ ), .Q(\u_reg.rf[14][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06622_ ), .Q(\u_reg.rf[14][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06622_ ), .Q(\u_reg.rf[14][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06622_ ), .Q(\u_reg.rf[14][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06622_ ), .Q(\u_reg.rf[14][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06622_ ), .Q(\u_reg.rf[14][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06622_ ), .Q(\u_reg.rf[14][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06622_ ), .Q(\u_reg.rf[14][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06622_ ), .Q(\u_reg.rf[14][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06622_ ), .Q(\u_reg.rf[14][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06622_ ), .Q(\u_reg.rf[14][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06622_ ), .Q(\u_reg.rf[14][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06622_ ), .Q(\u_reg.rf[14][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06622_ ), .Q(\u_reg.rf[14][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06622_ ), .Q(\u_reg.rf[14][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06622_ ), .Q(\u_reg.rf[14][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06622_ ), .Q(\u_reg.rf[14][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[14]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06622_ ), .Q(\u_reg.rf[14][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06621_ ), .Q(\u_reg.rf[15][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06621_ ), .Q(\u_reg.rf[15][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06621_ ), .Q(\u_reg.rf[15][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06621_ ), .Q(\u_reg.rf[15][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06621_ ), .Q(\u_reg.rf[15][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06621_ ), .Q(\u_reg.rf[15][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06621_ ), .Q(\u_reg.rf[15][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06621_ ), .Q(\u_reg.rf[15][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06621_ ), .Q(\u_reg.rf[15][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06621_ ), .Q(\u_reg.rf[15][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06621_ ), .Q(\u_reg.rf[15][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06621_ ), .Q(\u_reg.rf[15][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06621_ ), .Q(\u_reg.rf[15][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06621_ ), .Q(\u_reg.rf[15][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06621_ ), .Q(\u_reg.rf[15][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06621_ ), .Q(\u_reg.rf[15][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06621_ ), .Q(\u_reg.rf[15][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06621_ ), .Q(\u_reg.rf[15][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06621_ ), .Q(\u_reg.rf[15][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06621_ ), .Q(\u_reg.rf[15][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06621_ ), .Q(\u_reg.rf[15][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06621_ ), .Q(\u_reg.rf[15][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06621_ ), .Q(\u_reg.rf[15][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06621_ ), .Q(\u_reg.rf[15][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06621_ ), .Q(\u_reg.rf[15][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06621_ ), .Q(\u_reg.rf[15][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06621_ ), .Q(\u_reg.rf[15][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06621_ ), .Q(\u_reg.rf[15][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06621_ ), .Q(\u_reg.rf[15][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06621_ ), .Q(\u_reg.rf[15][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06621_ ), .Q(\u_reg.rf[15][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[15]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06621_ ), .Q(\u_reg.rf[15][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06620_ ), .Q(\u_reg.rf[1][31] ), .QN(_07628_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06620_ ), .Q(\u_reg.rf[1][30] ), .QN(_07629_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06620_ ), .Q(\u_reg.rf[1][21] ), .QN(_07630_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06620_ ), .Q(\u_reg.rf[1][20] ), .QN(_07631_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06620_ ), .Q(\u_reg.rf[1][19] ), .QN(_07632_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06620_ ), .Q(\u_reg.rf[1][18] ), .QN(_07633_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06620_ ), .Q(\u_reg.rf[1][17] ), .QN(_07634_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06620_ ), .Q(\u_reg.rf[1][16] ), .QN(_07635_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06620_ ), .Q(\u_reg.rf[1][15] ), .QN(_07636_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06620_ ), .Q(\u_reg.rf[1][14] ), .QN(_07637_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06620_ ), .Q(\u_reg.rf[1][13] ), .QN(_07638_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06620_ ), .Q(\u_reg.rf[1][12] ), .QN(_07639_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06620_ ), .Q(\u_reg.rf[1][29] ), .QN(_07640_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06620_ ), .Q(\u_reg.rf[1][11] ), .QN(_07641_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06620_ ), .Q(\u_reg.rf[1][10] ), .QN(_07642_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06620_ ), .Q(\u_reg.rf[1][9] ), .QN(_07643_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06620_ ), .Q(\u_reg.rf[1][8] ), .QN(_07644_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06620_ ), .Q(\u_reg.rf[1][7] ), .QN(_07645_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06620_ ), .Q(\u_reg.rf[1][6] ), .QN(_07646_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06620_ ), .Q(\u_reg.rf[1][5] ), .QN(_07647_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06620_ ), .Q(\u_reg.rf[1][4] ), .QN(_07648_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06620_ ), .Q(\u_reg.rf[1][3] ), .QN(_07649_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06620_ ), .Q(\u_reg.rf[1][2] ), .QN(_07650_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06620_ ), .Q(\u_reg.rf[1][28] ), .QN(_07651_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06620_ ), .Q(\u_reg.rf[1][1] ), .QN(_07652_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06620_ ), .Q(\u_reg.rf[1][0] ), .QN(_07653_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06620_ ), .Q(\u_reg.rf[1][27] ), .QN(_07654_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06620_ ), .Q(\u_reg.rf[1][26] ), .QN(_07655_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06620_ ), .Q(\u_reg.rf[1][25] ), .QN(_07656_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06620_ ), .Q(\u_reg.rf[1][24] ), .QN(_07657_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06620_ ), .Q(\u_reg.rf[1][23] ), .QN(_07658_ ) );
DFF_X1 \u_reg.rf[1]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06620_ ), .Q(\u_reg.rf[1][22] ), .QN(_07659_ ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06619_ ), .Q(\u_reg.rf[2][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06619_ ), .Q(\u_reg.rf[2][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06619_ ), .Q(\u_reg.rf[2][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06619_ ), .Q(\u_reg.rf[2][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06619_ ), .Q(\u_reg.rf[2][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06619_ ), .Q(\u_reg.rf[2][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06619_ ), .Q(\u_reg.rf[2][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06619_ ), .Q(\u_reg.rf[2][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06619_ ), .Q(\u_reg.rf[2][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06619_ ), .Q(\u_reg.rf[2][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06619_ ), .Q(\u_reg.rf[2][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06619_ ), .Q(\u_reg.rf[2][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06619_ ), .Q(\u_reg.rf[2][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06619_ ), .Q(\u_reg.rf[2][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06619_ ), .Q(\u_reg.rf[2][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06619_ ), .Q(\u_reg.rf[2][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06619_ ), .Q(\u_reg.rf[2][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06619_ ), .Q(\u_reg.rf[2][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06619_ ), .Q(\u_reg.rf[2][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06619_ ), .Q(\u_reg.rf[2][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06619_ ), .Q(\u_reg.rf[2][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06619_ ), .Q(\u_reg.rf[2][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06619_ ), .Q(\u_reg.rf[2][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06619_ ), .Q(\u_reg.rf[2][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06619_ ), .Q(\u_reg.rf[2][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06619_ ), .Q(\u_reg.rf[2][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06619_ ), .Q(\u_reg.rf[2][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06619_ ), .Q(\u_reg.rf[2][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06619_ ), .Q(\u_reg.rf[2][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06619_ ), .Q(\u_reg.rf[2][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06619_ ), .Q(\u_reg.rf[2][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[2]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06619_ ), .Q(\u_reg.rf[2][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06618_ ), .Q(\u_reg.rf[3][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06618_ ), .Q(\u_reg.rf[3][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06618_ ), .Q(\u_reg.rf[3][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06618_ ), .Q(\u_reg.rf[3][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06618_ ), .Q(\u_reg.rf[3][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06618_ ), .Q(\u_reg.rf[3][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06618_ ), .Q(\u_reg.rf[3][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06618_ ), .Q(\u_reg.rf[3][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06618_ ), .Q(\u_reg.rf[3][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06618_ ), .Q(\u_reg.rf[3][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06618_ ), .Q(\u_reg.rf[3][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06618_ ), .Q(\u_reg.rf[3][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06618_ ), .Q(\u_reg.rf[3][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06618_ ), .Q(\u_reg.rf[3][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06618_ ), .Q(\u_reg.rf[3][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06618_ ), .Q(\u_reg.rf[3][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06618_ ), .Q(\u_reg.rf[3][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06618_ ), .Q(\u_reg.rf[3][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06618_ ), .Q(\u_reg.rf[3][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06618_ ), .Q(\u_reg.rf[3][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06618_ ), .Q(\u_reg.rf[3][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06618_ ), .Q(\u_reg.rf[3][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06618_ ), .Q(\u_reg.rf[3][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06618_ ), .Q(\u_reg.rf[3][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06618_ ), .Q(\u_reg.rf[3][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06618_ ), .Q(\u_reg.rf[3][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06618_ ), .Q(\u_reg.rf[3][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06618_ ), .Q(\u_reg.rf[3][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06618_ ), .Q(\u_reg.rf[3][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06618_ ), .Q(\u_reg.rf[3][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06618_ ), .Q(\u_reg.rf[3][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[3]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06618_ ), .Q(\u_reg.rf[3][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06617_ ), .Q(\u_reg.rf[4][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06617_ ), .Q(\u_reg.rf[4][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06617_ ), .Q(\u_reg.rf[4][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06617_ ), .Q(\u_reg.rf[4][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06617_ ), .Q(\u_reg.rf[4][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06617_ ), .Q(\u_reg.rf[4][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06617_ ), .Q(\u_reg.rf[4][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06617_ ), .Q(\u_reg.rf[4][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06617_ ), .Q(\u_reg.rf[4][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06617_ ), .Q(\u_reg.rf[4][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06617_ ), .Q(\u_reg.rf[4][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06617_ ), .Q(\u_reg.rf[4][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06617_ ), .Q(\u_reg.rf[4][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06617_ ), .Q(\u_reg.rf[4][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06617_ ), .Q(\u_reg.rf[4][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06617_ ), .Q(\u_reg.rf[4][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06617_ ), .Q(\u_reg.rf[4][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06617_ ), .Q(\u_reg.rf[4][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06617_ ), .Q(\u_reg.rf[4][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06617_ ), .Q(\u_reg.rf[4][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06617_ ), .Q(\u_reg.rf[4][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06617_ ), .Q(\u_reg.rf[4][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06617_ ), .Q(\u_reg.rf[4][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06617_ ), .Q(\u_reg.rf[4][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06617_ ), .Q(\u_reg.rf[4][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06617_ ), .Q(\u_reg.rf[4][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06617_ ), .Q(\u_reg.rf[4][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06617_ ), .Q(\u_reg.rf[4][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06617_ ), .Q(\u_reg.rf[4][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06617_ ), .Q(\u_reg.rf[4][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06617_ ), .Q(\u_reg.rf[4][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[4]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06617_ ), .Q(\u_reg.rf[4][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06616_ ), .Q(\u_reg.rf[5][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06616_ ), .Q(\u_reg.rf[5][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06616_ ), .Q(\u_reg.rf[5][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06616_ ), .Q(\u_reg.rf[5][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06616_ ), .Q(\u_reg.rf[5][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06616_ ), .Q(\u_reg.rf[5][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06616_ ), .Q(\u_reg.rf[5][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06616_ ), .Q(\u_reg.rf[5][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06616_ ), .Q(\u_reg.rf[5][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06616_ ), .Q(\u_reg.rf[5][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06616_ ), .Q(\u_reg.rf[5][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06616_ ), .Q(\u_reg.rf[5][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06616_ ), .Q(\u_reg.rf[5][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06616_ ), .Q(\u_reg.rf[5][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06616_ ), .Q(\u_reg.rf[5][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06616_ ), .Q(\u_reg.rf[5][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06616_ ), .Q(\u_reg.rf[5][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06616_ ), .Q(\u_reg.rf[5][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06616_ ), .Q(\u_reg.rf[5][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06616_ ), .Q(\u_reg.rf[5][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06616_ ), .Q(\u_reg.rf[5][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06616_ ), .Q(\u_reg.rf[5][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06616_ ), .Q(\u_reg.rf[5][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06616_ ), .Q(\u_reg.rf[5][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06616_ ), .Q(\u_reg.rf[5][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06616_ ), .Q(\u_reg.rf[5][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06616_ ), .Q(\u_reg.rf[5][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06616_ ), .Q(\u_reg.rf[5][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06616_ ), .Q(\u_reg.rf[5][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06616_ ), .Q(\u_reg.rf[5][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06616_ ), .Q(\u_reg.rf[5][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[5]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06616_ ), .Q(\u_reg.rf[5][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06615_ ), .Q(\u_reg.rf[6][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06615_ ), .Q(\u_reg.rf[6][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06615_ ), .Q(\u_reg.rf[6][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06615_ ), .Q(\u_reg.rf[6][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06615_ ), .Q(\u_reg.rf[6][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06615_ ), .Q(\u_reg.rf[6][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06615_ ), .Q(\u_reg.rf[6][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06615_ ), .Q(\u_reg.rf[6][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06615_ ), .Q(\u_reg.rf[6][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06615_ ), .Q(\u_reg.rf[6][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06615_ ), .Q(\u_reg.rf[6][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06615_ ), .Q(\u_reg.rf[6][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06615_ ), .Q(\u_reg.rf[6][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06615_ ), .Q(\u_reg.rf[6][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06615_ ), .Q(\u_reg.rf[6][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06615_ ), .Q(\u_reg.rf[6][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06615_ ), .Q(\u_reg.rf[6][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06615_ ), .Q(\u_reg.rf[6][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06615_ ), .Q(\u_reg.rf[6][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06615_ ), .Q(\u_reg.rf[6][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06615_ ), .Q(\u_reg.rf[6][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06615_ ), .Q(\u_reg.rf[6][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06615_ ), .Q(\u_reg.rf[6][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06615_ ), .Q(\u_reg.rf[6][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06615_ ), .Q(\u_reg.rf[6][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06615_ ), .Q(\u_reg.rf[6][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06615_ ), .Q(\u_reg.rf[6][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06615_ ), .Q(\u_reg.rf[6][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06615_ ), .Q(\u_reg.rf[6][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06615_ ), .Q(\u_reg.rf[6][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06615_ ), .Q(\u_reg.rf[6][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[6]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06615_ ), .Q(\u_reg.rf[6][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06614_ ), .Q(\u_reg.rf[7][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06614_ ), .Q(\u_reg.rf[7][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06614_ ), .Q(\u_reg.rf[7][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06614_ ), .Q(\u_reg.rf[7][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06614_ ), .Q(\u_reg.rf[7][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06614_ ), .Q(\u_reg.rf[7][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06614_ ), .Q(\u_reg.rf[7][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06614_ ), .Q(\u_reg.rf[7][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06614_ ), .Q(\u_reg.rf[7][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06614_ ), .Q(\u_reg.rf[7][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06614_ ), .Q(\u_reg.rf[7][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06614_ ), .Q(\u_reg.rf[7][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06614_ ), .Q(\u_reg.rf[7][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06614_ ), .Q(\u_reg.rf[7][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06614_ ), .Q(\u_reg.rf[7][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06614_ ), .Q(\u_reg.rf[7][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06614_ ), .Q(\u_reg.rf[7][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06614_ ), .Q(\u_reg.rf[7][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06614_ ), .Q(\u_reg.rf[7][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06614_ ), .Q(\u_reg.rf[7][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06614_ ), .Q(\u_reg.rf[7][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06614_ ), .Q(\u_reg.rf[7][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06614_ ), .Q(\u_reg.rf[7][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06614_ ), .Q(\u_reg.rf[7][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06614_ ), .Q(\u_reg.rf[7][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06614_ ), .Q(\u_reg.rf[7][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06614_ ), .Q(\u_reg.rf[7][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06614_ ), .Q(\u_reg.rf[7][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06614_ ), .Q(\u_reg.rf[7][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06614_ ), .Q(\u_reg.rf[7][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06614_ ), .Q(\u_reg.rf[7][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[7]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06614_ ), .Q(\u_reg.rf[7][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06613_ ), .Q(\u_reg.rf[8][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06613_ ), .Q(\u_reg.rf[8][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06613_ ), .Q(\u_reg.rf[8][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06613_ ), .Q(\u_reg.rf[8][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06613_ ), .Q(\u_reg.rf[8][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06613_ ), .Q(\u_reg.rf[8][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06613_ ), .Q(\u_reg.rf[8][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06613_ ), .Q(\u_reg.rf[8][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06613_ ), .Q(\u_reg.rf[8][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06613_ ), .Q(\u_reg.rf[8][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06613_ ), .Q(\u_reg.rf[8][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06613_ ), .Q(\u_reg.rf[8][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06613_ ), .Q(\u_reg.rf[8][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06613_ ), .Q(\u_reg.rf[8][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06613_ ), .Q(\u_reg.rf[8][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06613_ ), .Q(\u_reg.rf[8][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06613_ ), .Q(\u_reg.rf[8][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06613_ ), .Q(\u_reg.rf[8][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06613_ ), .Q(\u_reg.rf[8][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06613_ ), .Q(\u_reg.rf[8][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06613_ ), .Q(\u_reg.rf[8][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06613_ ), .Q(\u_reg.rf[8][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06613_ ), .Q(\u_reg.rf[8][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06613_ ), .Q(\u_reg.rf[8][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06613_ ), .Q(\u_reg.rf[8][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06613_ ), .Q(\u_reg.rf[8][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06613_ ), .Q(\u_reg.rf[8][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06613_ ), .Q(\u_reg.rf[8][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06613_ ), .Q(\u_reg.rf[8][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06613_ ), .Q(\u_reg.rf[8][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06613_ ), .Q(\u_reg.rf[8][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[8]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06613_ ), .Q(\u_reg.rf[8][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q ( .D(\ar_data [31] ), .CK(_06612_ ), .Q(\u_reg.rf[9][31] ), .QN(\u_exu.rs2_$_NOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_1 ( .D(\ar_data [30] ), .CK(_06612_ ), .Q(\u_reg.rf[9][30] ), .QN(\u_exu.rs2_$_NOT__Y_1_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_10 ( .D(\ar_data [21] ), .CK(_06612_ ), .Q(\u_reg.rf[9][21] ), .QN(\u_exu.rs2_$_NOT__Y_10_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_11 ( .D(\ar_data [20] ), .CK(_06612_ ), .Q(\u_reg.rf[9][20] ), .QN(\u_exu.rs2_$_NOT__Y_11_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_12 ( .D(\ar_data [19] ), .CK(_06612_ ), .Q(\u_reg.rf[9][19] ), .QN(\u_exu.rs2_$_NOT__Y_12_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_13 ( .D(\ar_data [18] ), .CK(_06612_ ), .Q(\u_reg.rf[9][18] ), .QN(\u_exu.rs2_$_NOT__Y_13_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_14 ( .D(\ar_data [17] ), .CK(_06612_ ), .Q(\u_reg.rf[9][17] ), .QN(\u_exu.rs2_$_NOT__Y_14_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_15 ( .D(\ar_data [16] ), .CK(_06612_ ), .Q(\u_reg.rf[9][16] ), .QN(\u_exu.rs2_$_NOT__Y_15_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_16 ( .D(\ar_data [15] ), .CK(_06612_ ), .Q(\u_reg.rf[9][15] ), .QN(\u_exu.rs2_$_NOT__Y_16_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_17 ( .D(\ar_data [14] ), .CK(_06612_ ), .Q(\u_reg.rf[9][14] ), .QN(\u_exu.rs2_$_NOT__Y_17_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_18 ( .D(\ar_data [13] ), .CK(_06612_ ), .Q(\u_reg.rf[9][13] ), .QN(\u_exu.rs2_$_NOT__Y_18_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_19 ( .D(\ar_data [12] ), .CK(_06612_ ), .Q(\u_reg.rf[9][12] ), .QN(\u_exu.rs2_$_NOT__Y_19_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_2 ( .D(\ar_data [29] ), .CK(_06612_ ), .Q(\u_reg.rf[9][29] ), .QN(\u_exu.rs2_$_NOT__Y_2_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_20 ( .D(\ar_data [11] ), .CK(_06612_ ), .Q(\u_reg.rf[9][11] ), .QN(\u_exu.rs2_$_NOT__Y_20_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_21 ( .D(\ar_data [10] ), .CK(_06612_ ), .Q(\u_reg.rf[9][10] ), .QN(\u_exu.rs2_$_NOT__Y_21_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_22 ( .D(\ar_data [9] ), .CK(_06612_ ), .Q(\u_reg.rf[9][9] ), .QN(\u_exu.rs2_$_NOT__Y_22_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_23 ( .D(\ar_data [8] ), .CK(_06612_ ), .Q(\u_reg.rf[9][8] ), .QN(\u_exu.rs2_$_NOT__Y_23_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_24 ( .D(\ar_data [7] ), .CK(_06612_ ), .Q(\u_reg.rf[9][7] ), .QN(\u_exu.rs2_$_NOT__Y_24_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_25 ( .D(\ar_data [6] ), .CK(_06612_ ), .Q(\u_reg.rf[9][6] ), .QN(\u_exu.rs2_$_NOT__Y_25_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_26 ( .D(\ar_data [5] ), .CK(_06612_ ), .Q(\u_reg.rf[9][5] ), .QN(\u_exu.rs2_$_NOT__Y_26_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_27 ( .D(\ar_data [4] ), .CK(_06612_ ), .Q(\u_reg.rf[9][4] ), .QN(\u_exu.rs2_$_NOT__Y_27_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_28 ( .D(\ar_data [3] ), .CK(_06612_ ), .Q(\u_reg.rf[9][3] ), .QN(\u_exu.rs2_$_NOT__Y_28_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_29 ( .D(\ar_data [2] ), .CK(_06612_ ), .Q(\u_reg.rf[9][2] ), .QN(\u_exu.rs2_$_NOT__Y_29_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_3 ( .D(\ar_data [28] ), .CK(_06612_ ), .Q(\u_reg.rf[9][28] ), .QN(\u_exu.rs2_$_NOT__Y_3_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_30 ( .D(\ar_data [1] ), .CK(_06612_ ), .Q(\u_reg.rf[9][1] ), .QN(\u_exu.rs2_$_NOT__Y_30_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_31 ( .D(\ar_data [0] ), .CK(_06612_ ), .Q(\u_reg.rf[9][0] ), .QN(\u_exu.rs2_$_NOT__Y_31_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_4 ( .D(\ar_data [27] ), .CK(_06612_ ), .Q(\u_reg.rf[9][27] ), .QN(\u_exu.rs2_$_NOT__Y_4_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_5 ( .D(\ar_data [26] ), .CK(_06612_ ), .Q(\u_reg.rf[9][26] ), .QN(\u_exu.rs2_$_NOT__Y_5_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_6 ( .D(\ar_data [25] ), .CK(_06612_ ), .Q(\u_reg.rf[9][25] ), .QN(\u_exu.rs2_$_NOT__Y_6_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_7 ( .D(\ar_data [24] ), .CK(_06612_ ), .Q(\u_reg.rf[9][24] ), .QN(\u_exu.rs2_$_NOT__Y_7_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_8 ( .D(\ar_data [23] ), .CK(_06612_ ), .Q(\u_reg.rf[9][23] ), .QN(\u_exu.rs2_$_NOT__Y_8_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_reg.rf[9]_$_DFFE_PP__Q_9 ( .D(\ar_data [22] ), .CK(_06612_ ), .Q(\u_reg.rf[9][22] ), .QN(\u_exu.rs2_$_NOT__Y_9_A_$_ORNOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(ea_err ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\fc_addr [2] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\fc_addr [2] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\fc_addr [4] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\u_arbiter.rvalid ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\u_arbiter.rvalid ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\u_exu.alu_ctrl [0] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\u_exu.alu_p2 [0] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\u_exu.alu_p2 [0] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\u_exu.alu_p2 [1] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\u_exu.alu_p2 [1] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\u_exu.alu_p2 [2] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\u_exu.alu_p2 [2] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\u_exu.alu_p2 [3] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\u_exu.rd_$_MUX__Y_A_$_MUX__Y_B_$_XNOR__Y_A_$_MUX__A_Y_$_MUX__B_Y_$_XOR__A_Y_$_MUX__B_S_$_ANDNOT__Y_B_$_ANDNOT__B_A ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\u_idu.imm_auipc_lui [21] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\u_idu.imm_auipc_lui [21] ), .Z(fanout_net_21 ) );

endmodule
